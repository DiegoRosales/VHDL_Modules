XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��
�u�����h��������Ԫ7���[��7T��E���ߠU��2)Z����@$�l�υ��j�4D��)ҌۤfY�J�fg��_�T�ó ��r������\�n���i�(�s1n k���P5=��.��c�ys e<��ʭ/P��n}��]jDޠp�!�^�p����n��3xT���l��$ ���{&s�Q��^1��c�l4����-T�Ac"�u��A�C�	gE��3�>5ކNi*���ݰ�`�67;�r���_FX/y#��l���Ҙ[''d�~ӿ���uU���O���`޿�b�+��p$��r�غlFp�~J\�AT$ݘ�^��&]��K�*7IK�tc�ᜆ���͞���OcF���W�@��C%2�<��{�`>�I�F��m���ݹ(���*UpI��N΅�Q�0�&1+�|�0��?'�����F�E#8��J�=E��޸a���1�
�n��2�X�E��յV|LRG�承䀵���9�ۙ�`��&�� �m�+��X�*[�e+@/�[ڍ���IT�e<s�y/#]@.[֦�A�lh�l��BGGP�k�Ӥ)sS���y"��+�|�� �W�3�0��E�؝kzv]C�ER��i=�lN�_��N>�mQ�b.���gjeo�������՟�13�uM(��J����\FߔpŎ�t�w��W��L���@_��0T
����O����w��|�g�����ߜ��
�<ل�:oa|�*x��W��W��q2l�&XlxVHYEB    211c     b60�{�-P�0+�R���_?>~ ���3:m��+хL�[�a��f�]w�'K��W�Q�p�� ��#9��5�Y��+S�p�[���4Nw1�J��O�����C�����R��C"p^��a9ʹd�����g�F���7��-���s_`���{����Eh��N�F�1���LJ�a�.a�?ϜVʠ(�����^�S���<)\����2�H��KE�2j?Q+�t{�K<p�$��K)���7��c{��1BH9K�e��%%Bs���D�6��9�z�n�ј���#���x��7>yı��!�3��>y[j�GG�#w�_]�[����j���>J����_�o�)�ݜ,����S��8\'tX�QnY��6�!��[��������a�8�uaY�� ���7-�|�v�@UE��ֳ�-O� %�>h���#�k��_c}Ÿ�I �����yF�Qąp���*{B::���mz��$�ʗ�K���̆���� ��E埛}�C�֔7*�A�D VK�qN:^�X�A��g"�H}��Bʆ� X��`�92����Ϯ���J�7g��v58�N��F5F�|X{�P��W9�{������[Q=�	�F��Œ'�-���;j�e��$�<8t���e3�k��Y�M��nK%�A7�	.���'����M
U���������\��	��y�9y���ͮϘPϴSHD�5�xQ�2��Gn��A,�8��K4G����t�>�O�Sk������K3�#�,��9���͞,Bgi%��l��;7�?W6��x���s]�����atkj���빵S2��h�Ʀ �u͊'JS����l@��c�6�l<�Ki�V���p-|wX�`Q6>҈5��5c=V6S��c-�8I�U1�-:�{��*�2� ����I[�4�:����Ahc�?�����b]E���rT<v|ӧʂ�J���`�����U1�8��Pr:B��i�͐P:i\�r�kĠ���nTx�"�� �x��1���T��<�Z_����|���s��a*n����Q��XG�)u�H�:�!���`c�J!��P�C>��=�;���6�W��;!�!Z��8n:@ ������&p�d����~�^����p�c#��%#8��N�������s�l=\N��5�����G�,��W�=_�&�ؠ�e[/�BA,5���
K����ٻ[,��.�y���M6y���2aǋ��H����=@�g��݅)�Ȯ��-�D��������x���<8�y��$�dt@��	yfP�	���|$�>����枢���'M�)�+D���{����?jw�p�5�O0j�8kB����A���W"�= ��� ��z�ՠ�d�আ�⟛R��?6.��|5v���+�U�̩�BThS�Ւ��bm]����rX�?��3�n�V)\��+�����0ubg�����ڝ�g�'pO�\)�7��a�
��a�O��.Aݕ��&�g�E�Më"�??:�wY��<Y'(�O����Ei�4'ݡ=�~,���\y��`���i���׳���w6���3��3O�����P��S�������S�<j�\�M�6X9z3"�.�r��1m|Q�̴�Iq^�8�G��Wp�N�^]�>�|K�1Jo�DԺ�7⻰:�"N�������,~�"�b�d��m��a����ɧ��~o�V"�Gg(gTv�٪���;x����z��'E��E�g;��֦V~���,*��;��ڝ����}����c�~h ��ٸf���+��Z����"~㘇���g��������Yف���3RPӖF⣉!�?�T��#�y��$��@&�������YM)��4�F /S���L[�A%J����o���ks-OK�IC8�U��!��Ӄ�c��|�kG8�;��q���8C����b��t�\��:�M�m�Rl &�Z��`j�I}v�n��%�{s%�od��M#W�&-~�,���NVdmq�T4^��О>Q&��G�����#��|��}��v"t���<�͸�8woW�.��Nɉ��}+��ަS�K��V�C�B��zvLBѺ8LJ�p�9Щ��ˊ�/jz��l�={�I�V�F��؃���{!O���خB=�BϿ������n��N�:�_�[��{} J��f��t���^�55��(�����l�D���N�3�I�@[�]p��\�WQOH��I�+(R��{�=���������p��l�:�{��|̙Q�=�-�a���~���4&��qe�w*�z2��=�w��>͖���Q?ý�8m����Q`��z�uk���w�G������@9=�k&x�=���'��a����_ϸ��}�:�*3�/t��q��4�1��X�P!�����;�%�v@WD��ZIR��1��y9���2�d�D$�:."�kB{0���_%KWFow��%l�I%����-�o�_��Դ;	��X
E���E�c0����./��ə�,d��Ca�>*5*���A;��Rr�*��v(u��k��Ї8��q�o6t'}=�w���?b�_V\ǵ3M�� �Dܜ��q*pwI��'��0�)�ԥg�	@�Y]��z�5��5C�	Mz�J2�fP��?/���$ru��T�,�Ѫ�YςF�f�6
1�K����/oѴ���9�A�����n%-v��oS����q�9[�3w�t�����o��?�k�е(H?���~��������WCL�g���'��T7��
�2��Tې�??��N��F�N�s]c��=!�2ʤ�A��+��EEͷ�� ����/��5oF���N~�@\��71w	T���ۋ(yE�s�0���?UK�I�O��:��H��{����26�<�P