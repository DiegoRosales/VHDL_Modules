XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��|I�� �Ŭ�]4R&qc�b��_�e#o{&��c�����x��5- �/�P�ђ�i�^�<�o	)�8z1��e��4�^�&�wȏ�$8�E2}��(}g��]�Ŕה^��;X��u@�c�o֌��5����<��
*&�ad_�C#�؈�j�ߺ�yfW�_j�hͪ�+5��R��r�Mf�V��� Գ4�K�3�t��v�k�S�yHNA2��}��b�M4���N=��(�5�X'�!�q��kRq6:����:��[5ίp,���K�k��X6u&v�gޗ�2�6���	����
|d	s�]��� �T��.����&I6�Q��B@���Rb}��U�0_���)A�ܒ���F����6���A!����[Ҁ���+�D��\h�t�&!R-�u��kX��˚]�(]���$u@R�I�b.8�IY�
�!�엜d�X~�_"0<���֏���
F�g�#5�_�m㠈�,�?`sv0�ו��tJ~r��Xz�KU$(ԗ �ex�4'E�l���!��$����9���/!��Dk���3���a ��쉱�~���@[/.p�:K��}5S����z�!�#L��k��^ �V�����zMg��ң������7;/hӌ�����.q����&Q'h�z��r�fVw7q�>i=������/�s�!6x��R�$�6�g,��X�g$=SX�NްPP���1rU��ú��ʹQ��$�G,X��@�/��b>W���.���lXlxVHYEB    1ff3     b20�T�KJ�yjR�5��Q� �F(��W���ȔQ��>%��V�^�ɇ�\Zo�#^2��M	u1�k�)plU9�X|w��5�-F�g��S݂&H��BC�e��\�:����޿@>=���cیjJ��L�hé�G�
��?���/N�5�����{cw'Ni��
����C~*#�}�	���Um�#��}��[�(BS��0�����r�%�^C_����Q��?/�i��iI� ������
zLQ��$�Tڄ;f"�]<�Î[{\/�����w�̇�HR�*���
��a_���R�Շ�-�:������ĮM����t�>B^(|�N�:�m
���l���\7�MO����}��C�J�N˕��ј�-��H����!6p�`EU� pN�W�w��ZR��y!ȄDk6�<vI��s�j,���~{���ؗ��P\�73�~w�?�ev�S8��Ty��8��8�)g:�y��$r����g�Y��$Ŧ����?(�\����(7>G��^�"����T`R�+��/��(;��Mg藈��*�h.zd�%��f:[��b+���X��I�7yEߩ��zx�uT�`��/Y߮�D���(=���%�.GKϔ`��W�7Y #{���%�gN6���!�^wv��&L�PT,E�\�;��)�`6b�ڤ��j��y�p`z_���l�Oegj�6���zd�,�����Ƕ}��w
�<�[7����5�yS�͋-�[���X�_%��{�l�Z{-y�#Pcǯ�ۓL��)1P[���+���id���:��� ��� !}b a(���	���"u����N�O`/>ӭ>M
����4�����+���|h2n׶}RȢ'R)��w�@�7W;���z�P���-�$��Z ��R�����c��ǻ�N��|8{��X��%��mYd��8=����x�&~gH!7���CD�]!�������vaGj�ɿ�-/��G*�[��3�0�y���n����f9��<HY����N�a(P	)zr5�¬����k�����U��%5qRz<�zK��!a��w�kUd��]�*�95{��4[Dm�u���=.̺L��=��b�^
��ᴕ]Ի�d N�wr�1X��Ku��#�-1�u��-B����]�L�[� tk���}/WA�dv&�B�T�_��n[ct��~/��ǖ*�"�����=ZA����PJj����^�(Գ�y�e�uWVz�y���" ��V��X�Cl�D�>ʾ�N��üMPy�.p��u�Bmi�x��}$�W���~��0cl#Ƕ�ژq�}�å~R�mI ,r ��]�!��e��i|F�%�N�3�k������F�����5$ɂ]�� ���x<>e��ͩ«��w��+O| ��>�cJ�a0��Q���y���zH����F4�	��骄1hAC���/e�?3�,�f�;��S&K�7��#�ꑊv��n����Q����{�Lzj�=�u���d	[R��o��ۡ�|z�7��nq�6�����tfOD<���Zz�>�O8����M�a\b��w���	�{f����k�,Ν���e�Z,���G}����w�-&E��D����e�+�Q_�w�b!�/;�'��34E��r9�g����f�m9�I7�~�0�y&�Z�1	q%�Q���U�k��{W87g���E��;�*���Couʵw$�ym��_������eS�Lc66�(}�YJ����P.�����s�=�:/�[W �(�R�E���S�5!W��̊�3�D�{MH31�v[���Rb�c���7�'p�\(�vD��r+��
��k\g؉{rn�U�F~=.LԝȋۚX���V�[2�+���a��ٸ��L�R
�F屿�d��d�]O��Ґ�6�CP1|z:�� v;�� ��^����Js�b;��!+���Z\��"��쟬[(��5i`�x�xz~���+Y0��^�e�;9<�����G":���~�`Z X�Ζ��xO���5$��-��WJ��#0�[�1�@�� �jȂ�`���m���ꎆ+ix}���hѼ��m2���U_v��C5�_��AĴ���"�~�C:/^��C��E�����IX��8�G��q!�BJ�8�X�m@,�z��&!�8�I�ΚY:�g8��l��cf�lMGZ����ސ�����kNL���8��#g�\gʑ�%�:.����:l��+I��,FL������h�@ȵ�%�D�}���6#<~�K��s|���}W�Y�a:���A�1�9@W��1^[3@����&�E�GC���K���Rڐ\�!�_^]-wk�]i]h��4�6jSI��-�q��)e���8��e6( {J�R�1���ܳ5�NWۙ��)C���mע)���C�|�4�=��=p�v�r���w9��6�t�������n����K�Z�����P���@�� �DҔT'!\]ܝBfg�HB0�g�$H�8<��pfT%<����-�BF�X�#3v=�Ӳ}r��пr&3��6��|ϟ4�y5V�i��:���>I���ob�j���M��+�t�g3�O�ِ��/J�W���9燑tpvּ1�*�u��<M�_Ȓ���'���B�����z�F�f�d���,H�~����`Y�̩�Ҧ<����w�|��m��F���"#1{E�žE�����~L|&��d�g���8�����ʮ{b"{;!q�>�jkNX)���,~�h�$#�ۨ�E��I�v]�m*�F���Ң˯����4'(g��i7��cڳ	$&��u}W�U�4���O���Kv