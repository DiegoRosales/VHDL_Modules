XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�����~z\C"�ŀ6���$�1
�ef=�]��b2K�>��T
������n�hr�i�G�,�'^Ch��L,j%�s�fz2�jj��[�s�g�)"�f�����Vڶ֝�0�;��4H����ڀo�L���J��*=�H������n'n�_� W���k�b�I�A�%�O���vI�T�����2�:�9]T^q��rc����O�HA`Gf�5g����ر��!� D6}=�}nKIDg�m��株Ug{ۋ�
���e�\�A��U���HpPáV
�����q�MtE�^sv"�jT�J8;�$�q��k�H�M���n�o-��o0�����nq���=����V��f�:;��z��ݟ��s���c��^��C4)�nMkҽ#^�\Y��E���Q�d�1�X@n��%'���&��_�O�ɨ�- W��ҋhڝ���)��(jrM�����2�a��-��=7��DJ�F]�]�1��]���pLU1��(�2ܽ�q���#?�	|r���(�����$���8}���ާ��{Ɖ^����1�R��15��*�{r�,zOo��nL�35��8D
�{������\����tމW���@�J{��g�|7^�q���������`�R�xĩ����(�Uo��"��w�f��eCҲ�"T��01�!��"Cc}�F�*�]!?�O�~�|���u�iѲ�OT�Aoɞ�`d�,g�x��D�w#�f+���HMn��y�XlxVHYEB    1a04     940�p*�s��Ml�p��a���8/�HԼ��*���ْ�	��]|e��qع��Lμ��wD��vޝ�.éF�B��hֳ�$r(�<�"�գ�ެ�4����VF�BoYX���q?�٤�?����-,��C�s߾-h">�w3{o�)Tχ	6^<y��GOܡ�
ܗS�݌�D7��WlN�_^�`2����^K7�}*�u�R f��Ow�Ԯ��T���ؽF��e蹗�������D��\a��Z�	���j����tϖñ����>l�i�ތ'��Bj%V�.K����L3�X,�ɓ�� Q5�3ڒ��֓ �Hܥ�\� ���rx�ҿv!�{ܯ:)9�����y�B�EĂ<qEa���f���?ڷ�\Rv�D�W�q�-�A .��@҃�׈��2�O=�F�X|o�v�xh�\t�ӭ"-3�w���%F�g��|Y�1\�W��<�]������b���<��t=+�"iJ.�t������� ��[�Y�4	K���K	p��hz�2HzI4���i�=�^K��ǐ�ePp��L��g��y�~DTZ���`P%'(�`��,�g=�cq�s�$M0�;�x�B`v�]D+� g�Ϋo4�q�a����^Z�[��{N����B���E��YF�6"��>>vL�66�� ���+�$��?�}���ҩ�C͐C8%Y3�2b�qR�����X�	�/R�R�M��[��490�r?��)4��s�Tq��sB�1p��*�������6M"4�n	[-q\߶�`劫��;��C$��zr���l<	��|X%/�e��H����u8�0����X;�6�1�д�L�
��yc��%��yv�o_gu�S+���,k��{�C��=��X;8 ƾw�u����Z�0h;��G�i�gwv`���+��=9"�Hw8sb �\C�������"�c�u�:��_3��7P]D��p��{}�R,�ԣ)*�^�!�(KX���_�+^��I	��g-<au�X��ǯL����"���'#b��д����>�i!0����7��{�@<�f���-�#h��	^{l�������C����Ӵ]�nW��b��u��S1�!�^7�o��(���L�8p5��V)Rp�xD�����㬫F���l���{'�i(Otض�a�z���5^�i��OX���bJ����̔�!vtߵ�A(0�o��5w�cˉ����N(���K�_��z�QRl���ޣ҃��������,�%BnK�ؗ���"^��h}-M5e4�n�q,s�-c����WB��JI~mW�9���鏒@3���)C���~;IF�N����l�yӗ#t�d���7�61��us\κ~s��Й�Z'���E�QF���Fy�e��q�!S�}/�c��1�Y��[��d��N�i���Դ�2P�K���_�ɲ�zN�m d���d�R���&��Y}F�u�sP���P<PA (��Q//#oK �m�<�J2޷��8��6��.x�{�T١�b��K?���9��@�á�M(�n�b�\�B0��!]W�����TU���H�� �#!F,��4[�C�bfr��(-+Ā�~���p���(�W�$��c�<}nq�-�uhW�hm"�]���w���˶
�:%4�7�A-b�'���[_�۶u�TV�c�N�B��=x�E�w��m�zM�J�K��� ���E��9�K�e���������X�#$����2[�مQo_s�n(#����L�7Մ�{�k��}Nt���Q���|B<�C�g&]���&���Įa�64cs�!�'�+�Oj-� \�gp���ٮ����Q�|�w��Ɖ���[͍S~AԿ<i����Kdu���͞�>��#_+ڈ�G���$R�x5�VfC�Ўvn���@j�Q�!�8X��i} �-K�,oĂ|��IٟS�>�^�y�l+��R�~�t�Rt����1�h� ��$D���f�*]W�m}��"��b�+�;�;����.�����hT��շ]%w��Y�[��f��:�8џ�!l!+�7�#�X�0	b������:쿾cb���Z~i����o�r�*��8��?����;��g}a��Q�QP,��61�:8�Zy {�S4��F���(jy���}x�ŧj���چ����X�C��r$�4������b;�-�o�k(��ֳ���;��X)�8��+W�5嚷SwV�Y��.xW��,�;��;(�jTjc��
��ꅈO9����5�C���(�X�������� � aifBO�&Y?�E��ג