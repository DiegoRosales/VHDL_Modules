XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��͈5����� ��Y� �Y���ca�K�gN�ҧ���_
��*�4GJ�`#���<����a�R�#>��8��D�����P�#��$��5,�V𰠆���k�Y�>*Q-�(�"oQ�{�B*/�	���=x��}�H��K@�r=�[$�28�E�[���\v3j86�#f��XdZV����U�山-��5�Xl(�6��]	u�)��V⅚���$�7s�X�q�;A��G�5��W��t��������#��9U<a<�g�P��Fp�N5�a��C���mq~%�~3���u����- H+�C5���2�H�ݯ���}�W�r�C=���I�1�8&�t��Ꝫ4���)ߍ@��(����<��2�}�/����$�ܬ�F����I:�D�$RQ���C<�o��Ғ5}V�ʷ����P���q�Ӣ�o8KM��F(�|~��1^)�WɄ�y�F 1%[9�~܊z]��`i�W�t`h�^�+���p&*\����7/@$�� �b$b	ۢ��飰z�P:*vU4���K<��u�)����'^�6-�4AɄ��n��	�,W��ȦX��������n�C����$�zފ$��XW贿��H^�[�#I1.?0���!����սŇy�"J�U��A`��
����B���Iv�PNFZ�yᖠ"����V��Z�؅�{(�������c/�%�Kн�|<�D��
P��$ ����}
���t�^��4�nw0԰��XW��X��MI�cXlxVHYEB    2a18     bd0����Jv�=J������G}��j��ʁ�fՉ>�Z*���IS�h�h�O��W/W���Š�̊qZ��2w���B8g.o��`�N҃D���^���c�*^�׊p��G�,?�*�v8^A�<�d��X���}-��c���P���r���
ЅxS��e�g�����[EwI�%v��dzh预`&`�h��x]jw���8��#Ͻ��t��f�P�ؽG�+# t�s�#�.	X�#����lV�'����]��q��:!���\��Bf��Gj���|a�j�����7YRЀ �Y</hb�����etP���*d1���<�򞇞��Y��$Bil/x�VM��`�������N�ypu�E��V��B�N*)����Wdf�kN���73M��H���a(��=�ɬ~~k��,�ǽ�A��W2�% �D�q�T����$��@���b�n�$8��t��H{JS��SlV�*�x)�T�׸����B�"3�����x�ܹK��z�i=i6�؄��vH��QMu�}2�,,��R��6ї��cR��($+�o����.�@[����`�=N+�������b`��2s����<e�k�м6ց�VĐu�ơ���?�ܞ�t�lp
a���@���D9C��BNQӥ���z��0��ۣ���l(��i�Y¥,śD���Ⱐ���(	]���t�6�9H4�����^����X'�"�4p��!q|�ݡG0sn%�MFX�=��[���]�4�=�p�$�o?��]�0z��d�i�v!���x ��\ߊ��q˕3~�A����'\/i�����X���C�Q��c]��!n�I�6��X_ �q���LQ�:�R_\�`��QD�� vGd=)�����Z�u�6"�����k����G�lA�l�v������}h*s�ކ �mtB���ͻ�sN3�"&=�-��5�W������N�'Pi	���=.L&z-�YF��ꅷ.>�:��u�u+R� ��sO�o�(�++ �F�+��I�y�������	I��R��^���u�_Hl���(��|(�1#�����o(�ֳT����y�2u�]���k�֎9�{���=�B�d��>�����,C����VE�;0������d����IW_ 9RH�*p�X�Lc��*Q��~��O�p����]� NΕ�)A|E։��_e�9���a�G�&�c�gf�m�l�[Y^������*U� hŹ�Y�.�,��h��k�]�9%§'`��*ư��sV�i�NmOԷ��_Rtd̖��3�L���G���X�(�����|�
����t�k�XI��)l[����fQ�{��s�j�:�0ʀ>'����^S���xdR�Y�q���a�"6m-(,e�R����9XEԘa�M�c	�k�ͺ��8q@z�&L:]������Ӣ�
��P��[�p�L�ѕ�O�w�������t3Pz~a�I"�n�Y�'?�)2�J��]�I�Y�0��$֔����Y��+Y�Zw��3_��g"9���s8��L5S�H�.lX�u�1p �p�'��e�}����m�T;> �=�~��w^�&�db ������u3��Ķct�5X��R��ȋ���c
e<cc�2�aZp�n����]�Լ���S��k��=ڮ �ڙ@����ئYH�p�ߪt*7���H$�%k<6�x2�����1�R���̒�c&Mi?gfe'Z�ɿ��C��i�j�8�V�ۼ����ҡKC>�Z��թ��we�	S�I�	,�W�PƋ�Kw�Ec�I*k�9-�\=��iſ'���2j���F����i��M�������+`b�������j���P �*��,T����F��ʲ��=����.���G�B���΋ٜx_�no�xGS�=��� =�%�� J!��T��N����RR�}���bap��+������6��rz�@�A������"�)�/�{�����4����'&�#����� 6^�{}�(=#J���DoA�\��\�3�Ë��FE����|� =7�/5g(��IU���L���݊v;��aP!$�	�L�\�9�J�]Ҩ+�OT�N��џM�F@'x�'��HRZz@�NE�������ڴ�/E�rű-н�v��L�W���:V����fm��؎�i9���zA����,+
��-��*���Ub�B��N��D�����|���R�I=eY�g�[��y�p.����Y�{����+_��Q&)�4��>Fp����((�"*�\ ��g݈uT!�e�O�KM��=켋��ǔ�t��0<Y��G&rvH˳�{�0��3��M`�nǇ�>����8/6��)Xv�s�{���]�jr����1ޟx�+#b���FIеY
1*�g�j�
��ۭ��|�&��{e�$�C�˃�¾�JY�L<�n<UJ��#D-g�N�Da�Wm��}
��n�@1�]	�R�O:`�Y�>�����7��g+�a��Vs����l�Y9����z���&�8�jxzݎ��,b|���&��	;_��U��ی�4#s�6TH`9�B"e�� T���oܛ
[�F8�e�
�C[�5pxk�7zý�̣\��X�6��25�e�@�c|�#; �R�ZdɜwcڞQIhB4m�E�Ҿv[�B7ɚx��Ca"u`ё���$��$U+�8�S��|��略ǡ3���^�%�cb*3ঝ��h�uS�r n�����I#=���04��F�_u6e�n����,Ssko4������H���������C�z���ō`JguZ�Tb2�C!��e�L�r��@F��+����U��k��]GN��vo�o����:e{}1��Wמ�H���vmϵ`�29Q��mk����w q�<���y
��m�	ߴ��Oa"�����Y�k��@裇�����H-�����#G�(B58ސ�����JW�W�^'ɾ�5�:�y� �<g��twԭ�u�X