XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��<p&�,���-"��C��5jl�|�K}�?:��P�I^�k��� ��4�����4/��x�ї=��`��x��爥ؑ��X5��"�VU�a�1�%�I�o��)�&��O3e{��HA�z�> �����O�m���'j�R$sn����غ�� �P7�l���V��U��`.�ǩ��
22�tk�M���k � �qK�Y�T�B�n=���-�w���_j(���{"!hn��ᠫs&�n�
D-C`��b�h�mt�PI/��I�xU}���	���O����A�Q�� Ծ�ykK;/�9����U�W��wg�f0;dT�Bn�N�B�=Z��w����T�j1�qV��s�t���;şr��0@�2��͛;�����Ԯ�)��o�lrN��*h�e�U��Z��i�JT!� �U<��T����mCǌ^z�`P����8]b�z�q��$��1�f]1�-I�Ʃ�$Y^o�ejI��_��Y|�n�Z��
�
�i�/�L�
���]��ܹ[�*�'+HXɬ�|i⺣ìBd����L|��=�ދ��8�x�W��;�7�r�Ϗ�<�ڡ���^�A$��l[��= �"a\��$#`0�\��&��ڌ4ljK��)>��/"p%}?�H��k	P֛ރ/tL�o��D���徣����`9d�sF@�$Lpq. ��a���0�*i�t���@Og�ic �"�3�{�{VJ��pq'��Q�?>BK�������h��H'pw��}E��XlxVHYEB    5fe0    14803�v��X��A��?az�BЂ���ӑ[�3�}Z�pL�$~�c�1:rd�pX��im��_řI0U�A1?�ݿ�n*�DFQ�$�G�Q�z�J�Үm���|R��ͱ���|�m�� SE�d^���*١^aZ�4�����q֡��1�LJ�D�嵗��x8�i�Qg��9:����ȼ�V���~J���X׍sD��k���X�h� ���^� �8���|��2����qV� {���/��i2����֠�y3?��G��}�.�d�̚�C����ǿ\/���B8�ω��p):I�a\�zb�Pk�	
E�S�8����)��N���ʋ鐀���i�a��og3�Up��?�v�}W��$�93�%��|)m��vA��M���gl �9�,������Z�����h7�S��1TP�ȻA	��q�Ɋ��	����-7CJ�X�6X��S�#�O���|w� �7Nq9մ4��h� דּ�����n�ipt��|Ec�ŕ.�����.�HA`�'-�w���#@'c �)�?�5E�F�l@��m�&����_�����d8n�k�:7}�x���̪�:%��k
l^�yL؀�R����Q��W��5�=���{�C���D��@o�F�Lq�@����i_8��"�5]�Ĝ����R͎d��P.?\��&�'}k��:�Ӫ���.G���g�� ���K�^n;��{C!ߩ��X?<Y���xnN��%�c�Q#�E4�0�����������; ���2if���
�^W�3��������Rl#�W������5��ߧϥ�;�0�j�h��
S�mZ�c�U<��C�ؔ��+hmO²�7��!��K��rv�s�5�����(꼻"��c���8�����܄tұI�y
�k��,YPh�4�N�۵O"�+C�?�G�����q�ǛF�)G���O�!wF��t~͸����$Y-�.d�scD֊��ʮ��D:>��3�d�P��'�P��4���g�x�.8Җ��J�÷R��������.�ξ�	 ��i���J�=���Z"������[�;�q	EX"Lv9��	�}ÄL����2�J����.K߀{|�˅
`U�8�1�����N��1Z���Q#��KǠ���
=���N.#�!B*�%=�v�B�"�PK &�;E����G.��G`z���R2^g�h����L��7	Z�t�=5�xq��1m�������g�(��mû�\@{���o�o��v���:�D�	ͱ5��i�!3��Yp�mЪ����`�Z�,M�7�8&d��K��*�J��S^�O���+��7c���,:yF2�C_�D��G�5� �YnV��i�a_5��1Ʉ�k�z��݆o�?���"QW��=փ�35�d�����SC����ۚG�E���^��%A!�@��lq 29!@v(`�j�%��@x��:�&}<�P�"к_�P��NvT�����X|X�w�=b0��G���Z��t-�l�{��]��4z]�C5،��#�e���*Ӿ��N���QU�'�%��������g������x����˜��X��;���0<W���l�vs�5�T�y��F�J��~Z�ۼR��u�@�;�H�q�u�H.R�nTx����=zz��ۨ;^q9�Gk�2�t���%v����|��˅U�ۮo~�ӎ#( 4f��_�%X��j��M(�>W�ƌRr�q�pp��)���	��@�Uw��`G�u$�3��7���E������G�h��t��j��̠K�:�HD̮��� \κ�a��A�!&�Nt�Xe��z�� �D�:ة���]�+�3I1�����h��;q���F��ʕ	����t��òh�ԃ�/�U���>��*e�8{���HeI�~x�7��3�P���5��������9O"%[0�x5�2�H%���I�ȀlX �8�f�SR�a�{4�ag}�P��hFƭ��K��{j�����y���|���F�\�.�ue'g�``�u"�X�F+���4x�&����k?Ɋذ�6|C�Z�D�3
J��LzVm��^�_;���4��P�*�4bɩ�"$Dw�mx�� B�Z�́E��C8%K�^��B����l͓-�oy��Ufz���ё���1�Z�J��!���D�XhW%G�	|4.�%	[:�{֢z��P��U�܊y� @�����.�����*��i2���S����i��V��Z��hQ5<��ɛ�XCa�=���l,�ᄇ�I�Ծ��h|DU�Y5V�ﲖt�,���+�C�r���$��휹�k�L���X�a��)���\K��K��L�ш>�V^�t&��[�
�;�����ë��H<�cɽ�L� ��>���W=����!"!8J�w�0�f�³�[!1_������8�~�م�Z�5:�\]��Y��6���O��X��x]xR�r|�|pR4=)�S
�"�I�s��V��b޻����w˵�	EPrwiNG	cI�U��W�ͱ΢�mR�	RBKBO�M bn���sh5XI�+Ti���DMK���ޗ>���Hb@b�6(�F@�vD����N�3_�d����ӊ *�C���*��1�H�_�
�����	�w}���Q쫠�Ч�Y�:8V�(��U�}]j���Iu�hQ4�3t�%��pc�C����v�R?�m�s\�r�e����3%I�<�AU�]U$ބ��m�a{)70׶�X�U���Xڤ��؉��<gU�� ��NӉ}�F��D�|�1�w�:���O��(��tWmm����TҹwrT����J����s������e'�ӧ����zw��cN��f�����ӏ��'q�*�$��h!��6�$ol�֏��y���[��:��������nj��)m�:� ��{�t�R�?����܅����܉ɰ�曋�������{�����L�5ĺ9�il�pf�5��l��a��TEa��b&	�J,7>@�cxH;v�?�x���H ���xfS��9����8��=���%�7������c_
j|/����tT�|�ҳ��k
��T�h��q%��½ZFҀ�p�F��1&# ��{�T�K��աd��_�A��1H���'�DSs
u� ^�m_��&ƞ�h�U%���W����Y�TN�R�q1��]-b2�KQ�59�}�%�@Yη"F<��Ѿ6��r��i��p��S��s>bg�!��s[�]VR^ٔ�`d�������׌�4-Z�V�]�٘�P���3ߤ����n���u�.�QvW��Ɖ�X\��\���	oe���L2~�Sb��\�C� ��yǳ����[���nPӚ'M\��`�Q_�kg��&f�U���@��]3�"2$"|ǔļ�#}���(ޑA�u^�����g�(Lf۸L5/��
vÆ�kZ��X��\R҄M�Q����А���6O���W��Zl��Ls*�<�-&Rh����I+�0�c�'8׆<2o���T5)�?ߟ�_�e��u�K8�_��k[��ƀr!���������E�N\g����M]?���)5Ȫ�l����D�!.�dT���:�Q�jmu���Y-<?e��C:��� LK��,[>8���-��nnʕ�8�}�ǡ���q���4���IҢ�ꖸ�S�n�5D?�w��K'��S�j����
X|��@IaZ�0�Ǧ[���d��92�N+���ƊHjVWkT/� �l��ڧڢ��w[�����#�>���vZŁΌ�8��h=*`�}���qy��	�4]�?���^X�D`��\��!�"��,�>�qj�v�:=-��4;*����K���%|s�j{�I Q��f���D(eN�kd�5��޻*" �������ȩ;�=��na|V2�N
֓��b����F�'�U�nJ'w����>�g�{^mP��*�{�I��:��CI�?��&CZ/c7*v���o�:s/H��: QJr�k>3(���=EI*�7���J}��a[���nq�M�VX��׷��E �|V̉����j��>�Ț��g[��ծy�\l���cS�-�x���f�J<�th�@pI���Pش��o��I��*l�!6*�A���o
�e�U����؜,N����V@�]�7�|�r&9�l[��'s�J����;Ip/�8�v�K/��ЖLl���n��Qm)�)��ڽk���~3����}w/d�x%�=,���~�q���ڵAQ��Y��a�U�G���� �L;�ʃ�w���S���>��Ky����ضQ��z�F��ũ��9�s��;�����3����'l�=m��|�?��/�	�<
� �T�%�z־�g��w�O�a��=o%wf���0*�c��I�� �����to�1���r�ߊS�\Fx�+�K�S��H���7�-���x��<����z��8.[����.�ߌa��H���)"^"��qx��=���)��g�]�:5��1��l��xAzĉ�"��L1ؑf�`kf�e$�+a�sn`�e�Z����c�
>�i�·hNx������CH%��a��0�5����Jx8���g���&���"�_n�e�q��sQ� Ӟ���H�l^��ũ=c��j�򢲤����9T!g��$�L���� ��?
�6'�\�M�C��g��VZԛ���݌�V�|��d� �%�PF`�<�1x	*���w���P��
�'�FI�J�ϖx�oȎ���A�6MS�
s�]���#��6�XD
N�^��x�3&�����jl�����ߧ\�`�֥t]3kDs�׊�0bV��*�����V,F�Q�C��[����[ߎ�Y=C̱��BN/����5���;�,�e��	���[N���B���h��7<���b�L�e_���S[��:�ߖҟTF�vg#`B���)�W�,E�O���3�ri:�Ҿ@�������_��
�"�SF�Y)\�t�<������#��Կg�rCA�T��)(�h���I&p冺pg��J[v�~�2ru�*oFO�ml�[��dk�E[��ǿ7�x��b4��T+ݧ<�o�é�C,�:Ut�K�����ƪ�F��i�Ccz=����A��@����E*�ơ�� 0��zq����t���i9�D؎/:�����)Ni%�
�� �A