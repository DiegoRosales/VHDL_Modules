XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��cK�o���E����t�j�*����|$D���x瀅Ig�d��5��3m����+���>P��6��Ӕ9c��Il0�N������-���W���`�9���T��6D��S�d�P�m�kH�cO�	���O��v�16㝓W;3�0l"�I�����a��L�u��~���|����`_�v��|�GE�Eveb�e�/��Z��z4w2�!��{e�ky�j�i%/N	K�\?؆k���f�،B2u��I~�8s�+���;��}��C�nD�w/P�Y_lL��7�$��&���cD�TIl�L����4��V:w3�1~;q��A
-@}?���� �Nh�-��JBO�5�X\�U�#5M]����W����o�g�ؕg�24�j7ǈe�r��7�՗��H{2R����ڬ�g���a7��1\�N�-��H?��C�[��'HV����'Ãv�U䀅�9��ѕu*�T���C�7�a�"V"����+�-�d�?ɠ��ɾH@����V��Z�ᲠG�f���93v^B5"l�Ԙ�p�
�T̫�E����Y�&�r����g�/�<�Pu����X)�~��ɡ�A�h�R0�����u�ȕ�nR��j�XO��XǕ���ҋ#!���J+�δ¡���.H���}�����S��l�D73\̶ߏ��j�qHzHƜ s-����N����?�]��R��A�7��ui�OV7U��Y�0�lܞ�+�wx�H���	��U;�a_���!�{g�XlxVHYEB    12ea     7707<C�@�U�{�T��,�MaS�_���_�@�K#�//�i�֏�wj�}o���֭����|�fk"�j���8���y��C��3�o�y6'�b�å 
����U�}�=҉&���tב@�Vu��Ct}[�������*9��b[��#2���J��������F��|�a�:���X�n��9��a��ak~�r�A��=��t��6Y����c;�	���Utҝ�I�����UN ,�7����Ĵ�_�r�6�T���NR�*�?��2h�pJ�,#O<�m�_��X?�d��������>�����	������p
Q
#�0s~�H�<�����E>PF���;��o�ƛ=j+��%ls���*�-M�k���U_���dIs�п}�pa���x4��T,#�R-�vϓ����|r�;W�r�\���xv�0� ջ����,�����L�I!�� A�ю-0���59,X&hR��!�>r���P��
��yr	�D����_�*�:^>l�E@{ \L�������������49o��J(ʑ������XIO2�$z�r㋚�9�V588Xt�F���x3��?��R��+�}���@7#���R��^��׸K�"�&d�1��=K�\���{�^$@!2!������]������IH�n�B%V��S��Ѷ���[�'��=���E9`�2�^���$s����l�!I=t��������G��J�
>�D�*���7P�!�U�!i��?w/�55]�AJuǈԎ�e�9Gn1Rc7T,!V���"��CP[�>Og�_������ ���"#��%�&�Cu�P���2�0�M�41�G��̐�ʯ*R$��.�G�]���c!� :�(Oh;�H���ȱ�E�	z�˶�2ɽt>���_>P^���Zs�f3?��U:�笔]�2�4�
��ի���k%�$�8�:�����xD��) !�"a.�Hb��E��j�T�F�u��S�e����g�[d��-����Wc@eN޲��g�q��]L|ڣN%b^�*0�Z���K�v��69�E�;�%cw�7G�m�o��(�lǔC���{�H��\I$�n)�*t��D�ܫ*6a�����IYk�w�	������sO�bO��]�K��M
�3C,��!�K�4�=�>7҄����ޚ]�u�Y������H{i���J�F��8�xpG���7�3K�JljP���k$[�B����hO^�X[���$��o#O�	Y�V)��u��4�D2��'�zܜ�o����xg6r��8��*^d�����D�"��,J��,V��:��0j(���<�� �����k�{@�[�)	"�?��aF�G7UIZ�uc�!8���?�W�"I?��@�^eI�Z���}�`+)]�Nf9��)e���'�=�j��,�#|^\8KF\�r[2m�gO���J�y	
�5p��NmT�T���A�����7��Fx�R��./Т=�!�s�}���Oz�����s���h���F��P��-�h��ܾLE������%���OܳU�Ft@�$J���N��~ā�����策��b}7�e�\_?��]��;g6{kF�_[{��f��C������+�/��m�(��ߑL��-%4���fy޽����H�k�(��ԝA<��c#|<��7KM�f�˘OD�N��zdnA�b݈?]t&��Ý�mТ�&B<�oS8�� YE*�z0�ey�ݱH,���>�Mgh�	�����U�� �P�RL�h��i�%v1����;�c�֯�@�����>b\���yi�Q��L���>ȭ��.�%sn��vM�