package MC_25LC640A_TYPES is
	TYPE OPERATION IS (RD, WR, PAGEWR, WRDI, WREN, RDSR, WRSR, HOLD_ON, HOLD_OFF);
end MC_25LC640A_TYPES;