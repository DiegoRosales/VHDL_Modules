XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���gݘ2��C�d�u����5`�CW3��D�q�$ r7���Q�.���C"m��:u��� ->B�HD�Kӣ��ǒ-A�Ç<F�WD�<<5�D^ܪ�����)�;:&������Q$���ЛO�� f�ȃ�[F���>T���Tc4,�K�8������� ��v(!7�)Ce?lj�QF��}S�~��U˺S�}�^K���ID6��!7�S�F z��_�}��<:���B�L�,a��ke�؄�8RgT�KNF�����a.VP�
� _~D~�U��!��߇�Q��'�7n�2��cy����b�/�b�P�O� MIwuZ�� 0&�ǘ���l2�\���p�a`uK��f�mQ=W��츟��m���u�p
ս�dy�{�?��ӮAI<���uQ��Ю;�Ɉс:�`�3y���jRF���q�r��&yeV���%��>��f�F�w�VJǹ8����-�AuM$Zf�Ě�. �¹"�DhƃN0�F��%,�3*pDn�UHi�Q��Wqh�Zk���p��d	�G{H��[	�͒���y�ι���$H�8�b�sB�MW���� �i��Ϛ*G�OJ	�{3jMp~~*4�^��f0d;�B�=�g%��6�Nh�+2#LQ XӔG��45J~���O��F���[�`u�ZLmxu�n=qn�[:5���H�U�o�.�Q�q�<��2K
"���h5�9���zf�J���S��n��Mw�.�C��N��p��2XlxVHYEB    2ffc     d00��G�QwSz��ܯ5̘xvR�#�\�7��h˅a�mztK[�6�&�4�� òz��~@�{̦�15��0�F��OZ��j�>�����b�������ۜRຣ������Ħ[��)QǋwFց�}�%��*n$��޵����wz��?�e�.���0�Ѓ��XE�F
����:�� ���e`�����y��;��Yp�\쀘�<V��(^�^aP������e�8�� A�:��'��-28N�eL f��5�F\�#��$�e_�PD���m�L.���h�3���vn�� 7X��mĤ��t68���>Ǡ{d�F"D{cjc۽�H�WKa�Ã�mSn�\���L��
e��]�Fb���[ⵉ2�H+J߮�Ov5z69�4|n�x�|4���0�Km�I�خ"��r�:�!$܁&�^/�T֧�w	y��Y�����*F-�k9�{)�8����Ӭp.�c�����q���e@�v��1�Hy61�"	�?�ڳ"�!�l�)N��`
W�udŭ��:a��m2{4���)�=ěN6�^��#�Z%*��Z�F\�>I��H��A-���%������wV�o�=qf�Ym� �����5�B	fT+`�'z^�#)���?Q�-�Y�5�U��F)����z�������v��&�X!��l�&�� �R�Xߥ�g'2B�5���/J�.�g217�C�[ �1э��N~�U��b6j�Nh�����U������V�x�T������{��aY�Ha�.��a��A{�C�G\ �T�#m`
���k7��+6&s� �<�R��@�;���a�c1,�=�G3������a��4�8����w��.X_�dEF �bC>p�Eħ Fz����s��Y%�)::��7* 
.�N�#7���atg�(�HN�}N���	�50.�4"xm�����'j��i�ޜ����Y$M��ޜ���OmPu2zjhD9{sY���;��ښ^���Ϗ�Y�ƚ�$ǣχ'�z��g����W��6PS�v5�F�F�j�x,�������K���KX���G�����z�n{�$ޞS�Aa)�f�F�k�ҿY%#�Ei���]>��CA�q�Ň��>�fo�U��Ɣ�%���Ga}�o~%����O��D�*�:c:��t��0�!t+�؉An����QC񀂃�S��]�pũg��(Hʏ���n
 ����S�5� �!!,��8Ƣ+ �o���!��N����޲82�{MCAX�?��U�؏�{si-ޮ8G rXZ�?ocp�To��lZBe��� �>E� Y�u�Z˧Y|qhC�\ǆ���D#ƨ�ӺL��K��6��/�fȰK��9ER�[�EF�<>�J�ܱ��>�T3�ME�5�Dt�&��:�h�i؜{��c����<TnNB����)�Z������X}� �G��9��`�|�^�0�胭��J������\��D���g&.�EnssI_$MN�$�7��7��yZ��=�"�Єw@]�s}��S�f�ճ�U��O�$s_�=):_��A�/�G�}#�HS����_��&~2zM�@�	����ӷ��U<$L4!��'������RcųxS�P���u>��Xu�e/���P�^�+<�<\\�D�{%����N2�1��A�A�ߤ����\~vw�������R������m�ͺ��G�f�78~s��6J�	qۙ��^�WțA�U>ʗ�;2;72ޝ���Y�P���̈v2�Rڔp.�xXi��du�4��E����C�*E���ɘ��{��z�z	��|�!H���$�������ܵ�.�@ +��Bq����H��-�_|��if�K�:�.l�������C'�N<�q�R�e����"�-� ���_� �	��䂪&	���*��p��*�9��������M��2�﯅cV��E�	Ѧ6	�3����~����'�,_��h��v�;��D�?��F�Ñ�g�a�<}ރՕ��@!cPRb��ڡH p��1V	"pDَ�|�+.� _}���
/���Q�B�Hѫ��4��JY��wW���"C0����Ұ��D,:Bv���|l���A�)�5g�{��ş�j�K��,�|�g>��AY�ᆪ��42�P�����sU�Fω
}���{�l�M� -U�󜱯k����I����a}���Bc�I���Ϲu�b�":��s�K5�L ]����r�P�n��i4 �E����d��� ��۽=y��Ԅ޻]�q��M���Fp��E|�K'w�-�$(�N���\l�����܍u��e����&H�}�1��bY5���l==
	k����D 7$���&�����3#��w�����ؤ���=�!R8����l�0U�2꫽s�*M���IP�`���Em�[���J,��0kA&H��Sd��"��A�Wi�Co�� �Y�_(u�D�U����y�8�H�E�?OD+=�/��Gz��qu.R7ښw,�E��j�SX���[|�<z
.U&��0�R���E�nc�rk[�f=�[N�`i=u��)p�ĥљlBL5�d�k��#m�Zi=7~��@�Kq� (0���\�uɚP�M�p��W�e��������g��5������}�cn/�I�$�j��o��lܵK�\�����Z)<��wX�y�b�CZ�� �U��˝�/�<�e<�N��9�XL���T���Ny��~a�d��|��X_���p'�� ,����3���;�<��8Be��\I�Y�`�И���͸Nb��"�b_Ǝ��2V���JQ��M(����Bߴ�!L��Ri��%45x���Ć[����J#�`HJ�;���!x�~#�AM�h��\�U3Ò�0���TD*��RW���n�\{��H�3�΍}�F϶���M4����HOMm�)]8��WS�ݵ�C!�)�s/rW������q/#��E/F�kF<t�>_�]�6�"J�D��f��U(1��릑��0H���v�.˪���_]E�w���&B<$D(˺���P=�W�b�W�b����7<��}yc�[��;R��+���Y�y�}�by",�'~i�/-pK� lA?. Z[��Z_d�Mr�!���.L�ۗ�9�A4�>yG2�ye�y��d��W�| ��_�܈U(����|�b�)�B�y�[��y(e���:7��'��ᄚk�p����6�o���4�pO���
o�N���.8ȿ