XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���������Z�
8�(}�<��^x�flZBx�#�;]�
W�c ��:N�s����t�����Z����*��ZH�G�2��o�]8Z��=2���??��bQ��:�l�+d49��C�����>K3�Vx��������(����BV�{���׀���cP�j"�Ĺ�dbi���3*�_��n��n�Y��k���=���족 6�����-���eġ�2�u�m�<ibF���'��ykF��˙F�����@�
5pl�A=��1f}*/7�#o�-P;��.���ˁ��{�=|h{�%�+��k�b��ޫS��Rx�'��*w@�D/X5���h:?�⽚7�S[S
�Nrz���4�Ds���q�+*��`A��(��2��I�������f�~��6�=�U�S�s��q�s.>���D՝����$�!�,�`5���ܱY�0�I��,	~PX�p╘C!gr���	t���%j(��88E�/�濖����)�?�X3�(���ZNlx��@�~���M���2L��'�;�H���P��Z=�ӡ�.g,a�Za�=��FܴߤV^o ��y$׹L�Qq�ڴ)�<��n���ε[S����6��ݍ�ss����MX/)s�w�( �Z[\��b��$;���Ω1�ݻ�i���Wh�V��@��_U���MO�Yh��I3�R����$írC��QG��48�����Õs6k���4����H����j�GZ�R�k�Pj�XlxVHYEB    3ad2     ed0��%�*�	�DO���xoeWf���g�ٳAZd¬
u`��|�{=��*2���:�~�3m9���M-��)H��;_�E��f g�?��K8�����g	�N˦�i����?��?i�j3��q�_�J���J�;��t�e�z��w	�~�����Vi&Po�/�_U�����P������������[Z<Ob�ܕ�%n'�K���U� #%_�������
���"mg��G�7�0�.��?�R��iyr�;n)	�gŚ��E�U���~A�7���M%��4�5� c�?�I��D�	�Nh�Jx�CK[��(�>wes	8�'��,�����[�
��Q&��[�&�~(MEd7�d����#���,m�򖭙��7��ڲ)�;�/�Y�t����*6|��@���|j��h��z��}o�_�����YQ��95�f;�FZ�tg�e��� r}i��)��:iN�A���d)���H��w��<�&ҫ����4h���&h�	����Wi�b��*z�f�2"b��sw4G��ֱt��g>�fG���L�I��?��_�(�Qi�᳎�$_C�J�!9_�
m��RVs$������!q�X�a�k+���� �e5@E0�R��ԉ<�W�"|�9@a�*F�3쥎�����F`�E��1�X�C;؊E�|]�_p��tF��}�}�5���7.�R�J^3�b��#�2�W�]l$Y�/��`�e\=m�j��Km�D��lq��_����U���d� ��7�M�Z@_�r��
Fc��*X�{���L��G�%v��4k|���_�%4f�-��wq����K�ꉨ��'��D��	��@�+ �\lbg��O糝�;2�TYwi<X��ε��27/�	�#2�^�A(f�p��Jg7�Sf��Õi���ѣfZ�7�F�0)��Aަ.Q�$U�	��b*�(J���j�;;S$(�AJ����;���ș�G�z{I-�J5���\����Uad] ��E����'ÝV�	QF�~%�X1&�x\�BS����h�n`hx��a�9�[�s]mBdAC�m���6�i���T��/V��8H5J���[�f�	��5�lBzc�����s����F���j��g�Zt.h�	�
s�]������=�f���H��+0��2�Ձ���E����W�N���#��+5����k��������^�A��H���^�sѩ����⣷E@��It�#�~���Ñu	��]I��A�=�Us�Y�9��}D�82Wv���5fŰ���|QW��ہc�C瑷-�����ガp��'i]3��b*G�:����	�p��^���tc�˨�f�-�w{k�r���N�%=C�n��:���:��� ���z��20����	�XɊ!�w�9�I����S5��^�;$C*d��[	�}U��8r�2sN{<�Ѯ�c�L�ჟ�"y�&�YUsGAl���{�r���>�r<�ߔ23��Z#ŰF^��$�:��~���ʮ������)����l��H�&�R��� ���9�1hvOB�A�CU/����6�@�
���a����xF zC���p�ŕu[L~�9�C*�Xҩ �N�<��"զ�*]�4�Ȃ�\pj�↧X��v�g"1���%4[kdVm�����.���9�
d����늋��sFv�
j�-��I9j���f��Ť2�ϣ�)i���S��z�L�\�EgCH0���)�b��R�/mb����N"�0�'�HF;�b��vU�Y8�	}b�V�~v®5�-@Og���]�K3$]����X��M�W9�h.��8��2T���]�o�^�$3�ȼ����7�H�i1�+�:'���mT��0�<@L�c�]���O��o��9�k�%������2U��1�& �k7���z8^Ð����fé���)U_��B���?B�,sի��g��{�N8z2d,���	��FZST"Q?�\HIZ�Fu��F�[���	��Yp���(�4�B(	C ��oۂ�� l����a��+û=��S���;I��{[�#J-��h��hX�wR%x7�d2X�����:���V/���B��cjF$�%dg�����.���{C�@X�T��,�U�f���'dYQ���L6�w_7� I��.�%��u��{;�-��z)��"x.�P ��:]��e�%O&�iOD(�%3)%�#�m���hrd����U�!�O�|������@�����7�v��<�������#��N©�?��G�K+�/TҲq@�Ÿ�:�G�����C�6i�u+b o�*�kN��*]�`&؆�&�KŨZ�&��<��R6�4 ]�cZ�|b��fXw��P��n���&t�gqh+�&�u���#"�4��(Y]���g��j����ſ�|�>F��F�$'����j�35q�eww�$�'?gq+H5|��""�|3:�>?��A0��u�.)pv,�d���%ȂyŤ��	1��	�qS�,V�oFQ��HGc$�;��%�?z'��Ct���saMv���0OĴ��١��b�/����Þ�������`��Γ1�C�x����e�|�/����Dĩ���_�;ך�o	�	J^���ԭ#l ��A�L��A��`@���}�](N7 �� }�+��HЊס�-/��B�b^zoV��oLd;�=(�?�R
(��{�텿[���[���QC�`�'������j��N�mA�L��4�ݴ@ܛ�G�񰋩>"����KJ���`�����=��&��^����/l�$i(��ASۑ�
u�M���L�ߔE�� ��m��V��Ԓ&������z�oܚA,(=$M��G��3�>gGA(C��0ʫf�s('�v�x]p3G��b߷���H����<�Jɫ����b��a�5Ї=�W��~��O��K�W�^��K$��ܴ�I|�{-\�㥞fv�@HΠ(X$��m�<������{��S���z}� IVu�_�>��xӕ��EE��G�N	�w�^���� N8�|(e�?,9��J�'�F����1U]���o$�l��]�
�t5HB�7��Q8�8�$D��"6�_�)�"�B�5C������%Y@�)�1A:F�\>4Ȱ,�������B��މ0�1�O��aV��JO�{PZT��1��֊V$��M�*Ω��@�~���Mc��k*�zh�em�0�K0��J!2e���AYϡd���g .�:7���SZ��F�V�yÿ��;Z���ё|���~���x��P�kuh5�j��I�⹛��&�M��s#����S*P���1z�5��
 ��LF�k#�H���R���ُ����!�5i���@^O�^gŁ��)����q������ 3ak	+�'џ2%�y���@5��6읩�,���Ŝ�s՛o;nT?B�;���|�����1q`�AY�;!�w���n[j�7Ñzd�FP�Q4��*��t���櫋ʽD�����r!k�}(����+����ڄ`O����;EgDѰ3!r��,���_�^е�g_%���DԎ�kH����c�q�W�z�o�X��*����~4�A3��̂ի���\_EwPز(�.r8����W	ƃ�H�hϨް�� f�1N|tX��h����z�����@���o�