XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��u��a�4��[#����o.v�Me�������0���Q�N�V>�I��I��O����$��j�i�ƱP}�}�%�j~�1�eq�T��<?�J��<� ��T��{��59r�c�:��/zOSd��D�����?���6M��Z�3pKǍ�A¹[F���+8ΠD��_��o�]��C-(�_6+���A[��
��ҸP��7��x�ϴ/�}o��LE���Ñp���!-���s����9:���q��K���*"S9�� ��Ƽ|�:���6�Ù�M���� �B�)eu�?�����7?5D˃����}�Qjضo�P|s�=L�ʩ��4�o�;�稑*�b��$[Ԍ����2�:��?�Z�Yw�ݠ%^����n�:� $?(w3N����\8ǳ'}�.��
�T|�U�Wl|f���g�T�R�>cC��8��
���8�,��7��ﯓ�-��|�����%5��G�)����4\�KTM�kQ��p�!x�Hp�
PC�������1	
�׀AM)N wx�7���r9|��&�U����5��K���ZЖ��S�1l�f#0��Z#r߃��I�����"���g�-{l�FV_���q�9��RwҔ�H�(ii	�C��u�&�ː����!|�7�22�4֍��l
��&:�{��I��W����t�3��N��ю���~Mٛ1j�{�B�݈c�B��%�B��լ��;T�'�_y��q�:U�p��	2t8��Y�M�XlxVHYEB    3c1e     f10������|�ml"!�u����'��j]� ���(,t>,��\�Ź]���wi�>��x�L��Ea<�f|[s���suh��BNY|���dj3�eK�ܨ���:�2��۫���MW<^{[����˧ 7��H���UJ�-*'x�K��Pf�h�4%��E<��o���G�}G���gE�|O��S�'�aՍ��sn�c������h<����b�6b�����<���a��;�,�_F��C���?����,��s����r ��S���x�mn��g�+�('�=�I	V?G8AЂU��:fGe�XRE�W�m�/T3A���,4��ro̲�T��p����n!�����ɜn�/��{�>!�$���yfq�H���B!*��f��*9��h�'m�>�oG����5�K�\ك}�T�.�Y�펌�R؄��m.9�c�����B3���XRE����ڲ���7���n6:s�.�{!*?�L��4�WD�@m�Fio�c�fNq	��J��|R�4�
��Lۊ�[#pM�Kє�+�J��hcߺ1�}�>�-�N�%�UD�{e<W���n��s!��'.;��8�D��+�Tly���UB8�B/M䲚"�O��\x@���g��mĨ��R�FƦԍ�DF-#��P!��:rs֔�����ɫ�Z�kC�77U
|��W�����7��=9��d1�LD����r���L�����6�m�4��&8�6��c ��0�َC�k��?lz`}^bj@�y�������M-�1"��]K9#�grLV,a�,�N2e/2�R^C� _�\6(�}���t�)�f��+����������FC�;c�ba?7{��ՙ�~�p*��G�ً��q\�gҏ.��W%(���ĞX�$��G�AHϭi��O��p��i�[Ұd]*f�`����GU�ˌg��O���E�н�#c��(:��c7��E^|��$�hG�X��be����u̎�������1۶�%�s��m�]�{7�Vj�[PHv���9B@G�������6=�\x�M\ׯ�A�5�02qh��a#�ז>|��pS�ɀ8����~�����S��A���n�p�	\�i�$T�>�
N �<�I;�Ы�n���#���/a���կc桁*�|{�q �8E�%���P��62{��|�"$�P/'""���%#��b���I�	�A��aV��m0R��.9�	nw���-4��y:x�Q6QC�:?���@�SeQ���q��Ҡz
�W}���b%>�ǫ�ӓ�j�b�.��G���X�#��	����ͫ�ŅTG�]|� G�)��1�C']�Bw`���D���	��H�Ҙ,Z-�̾�m'��ݒ���NĳOB\a��:�ab�aF�z����l�Xe)��Ps����aN&L`cU7:-��IB����2��A�5����W�̊�t䶺n�xv'S�K�sg7S����X�kg��d����~�OjQ"�����kRGi�<ө�\J7� �����iж�E 0؝�JxK�!D;ҴP$`�v����9��}�C��2P�(�T!wx�*�c�w����I��"�imi�y��r��� ��"K_��u��ѯ�'Mh�Čcl����Eiُ��4I�3�P۷��������c=I_�n�\�&�Σ�.N�1� e$`�Z��N|ߑ��`�P���U(>D(���S�&��'�Qw:ie�q����
�WHJ����W�	%bW��o���H#@�Ut�zM��o�w����@N^rS�L�O��h���,���,c�i��o��]d9����[^j�ի�O�o;0������-�t�LSJjm���a��iM���j�[9Mx.tn��K!ءv��4�k6��S\a>�������u�*�����^3hj[���E��N�^��y�!/��Ԛ���UP��ʏ�o��1-%���b���s����:�)/�N��,ΐ���l9�Q�I�T�$
��9f�Զ� �ĥխ}�4���š��\�.�*KD�AҠ�x�±�rґN5���T�a���F�9��]K[��2A~�ȑD�1��7�Ұ*)�Q�~��b䲻��cXY��:U")���a��K!�oz�qeY��	L8Y���|$���������b� u�E&P��p�x_��wb�<W`+���>f��_xcd���C�����tb6��е��_��6�[@����ۧeVj���� $�N�z
�<�k�I{��hS�q�S<�y�p���N�g󸔥�}�ɭ\]�{�iX�D��Wvs�	�>vt���SW/�j�
��I�f��ʿ�;��r�t�~� �3��t��eGq�[��+6&��5�8/L�]���^Mފ�]�*�P���|�4UĻKm;�Nͼ�$ݯC���ʯ�7o�����znk,�R�t%�6a]��2��t��t}ByM:���u�����k�,V8��8Ԝ�vm�c��ʇ�I
b���<�{(�_�A���Z<�֯a�ZC{<����Xt�wY��k^iX�vCl�GC�X�A���~�'��L ��f#1�&��<d�HrdY*W$��m �M0�(/����������L:9w����~=��nk�̈́��$Pt��zkP�$n��?�S�5@�wz���}�c9i��=g�c��9Sx/�ܒ�s���}��ɠ7��:�P�X��1���ԽȣM��?Olx�럈wIy��q-�s�e3QK�E�Ő���u.�s���X���ٱ0�ۡ�~d1tV'?S��*��X o���k��V�����n�q���P���T�D<�V���4y!$�_�z�L!�_�Ө����� &�/�������k�S:FpA�S�t�O�l���@�^�O(���|_T���Ĕ�����|&c�A���5εmj�����%`�[������lY�B�
��ˑ\5���h?k;|�M蛂,Wv3��
U�iN�l��!���a�� �:ه�<&��A[�K��}�rc�
)�3����N���U�`[�Fs%����*8� ˠ��K���4��N�Ǣ2X/� K+dLqu6�����,ApB�V�c�<SC�=5��vź���r���C�U���Î�^ح*ٲ2Eί�PA#iXq/�P8tp\�dL~�*F�E��bk���@,�r�̝�iLY؅�R~�^^_��(�je�����!�6$�3�Zz��#���0��#L��{���q�yvOC��,Ou�9|�,։��Ӊ6}!S�"��s���#=e$�o}��/[��<��f�����% D�.�����QxY�y�.���%�u�®�������9�J ���{M�s��;���d��t��f�8K��k���ղU��@f�tz�Y#��>8 �mNL����Z5{b��j[�|���y���l��ǜ>��`�YF��"�u9�n-3�F��� �5,�����S���m^ �2M��u�4b/�*U���Y����R4�����l��-�b(J���������aAz&5��� Rϡ���j�Y]
��CHKAJUk)��4#�oC��,!�)z10���H��!p����P�ͻ�'�,Vsu`�Q��ҥ�`7[_����8��XPanN��4����1���Ō���ɻzrE�*�+Iy����G�%������c�i�n'��%˺�l����m��_"��ɥ�f	`�㷯�m�VYV�G_���%� ��k�䇵H"�@ol~���ɦ��Ki��l7E8�H)7o�Π�&{�:������	C���XP5