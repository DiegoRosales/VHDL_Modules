XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��Rs�z���"�O���nx�\.���N�܏�q�(nd��/���Yg%�;yI��'�E���� A+�ɸ���Bʬ���0��H����7#l�˗Ձu&����W���9MH<</�����!8[�����a͗��<��-ua�>V��R�e��/��wg#X˳5a�iu�?��/�t'i�@������qd_�]�,�7K"�}m�F�4��!k&��#�A�&�?�>re�:H��{�Zp�mi�>� �����oM��mlL՛:�GUX�����kt���7�����\u�qr��N���0Zm~�W���x�N�S���������H��Z�0�s[�9KūLȶ��UsS���^�z�B��ˋ[��=�i
�p�1k�Y� 1��T�k�+��_����F,7� ���bJ���	B!��ˈ��pS|?I�G"�ڭ�Hz�ǻ+o�&y�����¨�+�s��"2��5̇�)?3.�� ����-Fhk�3�R�Y���z��1�8<���t-A��i)tȸ@�~]�wtf>������ׄ�QX�s�;�W�0ML�����biuJ�a�Nԝ�=׈�j��ɑ�)D�DJ ��:�@�x�R��H��� 兎 Н�6:Z�%�8�Z d��Ͼ���>�)Ν� ���k�AYj�/l?D��\w�'qd����u}2#B�2\(����0rP�zV;�XǼT���M�W�`Q���ڲ��c��f��1����;�5�1T�msj[,�XlxVHYEB    516c    1400�Փ�)2�^"F���p�wLU�g�r��dJ��:�(�G��F��>Z�l��yl�nlla��f��uY��CdK!8�V�˙�Af��~��	=�,�#���̃dvq�x�78��"�J��J�
dS�G�Nni6Pa$��
c&���vȍ��_K���'	_9,zߴ��F�jvϚ�R�īc /^/��`	ZQ��~���� �&ME�*��G���e���#��F����:5)��|�U�,$D��?/��QY��N� ����!��*��c($-ǻ����Eb�$J�ˎ�k�<�1�C�4ړ�إѓ?�D���N՘��J��5��T����"* �S�/��k��Nߎ3��	:�����>���-���+�-�g�v�2`��7Z��W. ADڢ��	�n:�ie��d9��	w�&	#w��M���7���@^�iTK�rE&�ɉՊ�/
ɡ��)��fp�O�>j��<���i`��m�ϛɡsv�	o�e�!�&_l/_��Wl ��B�WHr���P�Q��ӫ��4���vќ ��/�:^�p$��z
@�6���ˋP�c�N6+��gR�>�/�ss+����8*�'��m:�ϱ˕��)���+-uq�I��\C��(���qg�c���q(�f�(Z���bWK�j�����
;�GD�S_�o��&[/���V�u+�$��]�їr�������.��HSns��&5�>%��Q��L���j��_b"�'����Z�'�o�V^3 ��&�V�ji�����Q�AJ�- ��>��Yu�C!o⇫�
���*&�VP5zV�c����c�����N9&����g��D����vZ�դlk3���@pC�?�@��\�m^�wf���iK*� ��r�k��LC<��\h.�T,pk��9Q����a#v�:PT�c�}?) �LN$4r�����hC��M�C-�ਜ�_�r�` ��wxṰ<"1��9lr%
<�,* r>����l��&��rwס��7������t-�����]��a�Ī|J6F0f�j��
$�r�-��][��4��$i�vS�pfJ��7�󖯍�ECz��+�.;V�[��٩��O���d�D�2.��l��%V��Π�`�����q�IP��� ����ɾ�=|D��rݴ;ps�o5�E���8��w?�l2a*�m��_�Eom��i�E:X��HC9���"�P �^�������4��%���&p�nyzL�ֲN7��ӣ3�CB�2�7E$/�l��hE��a�k����d:���z�y���n���k��S�\�����#�)�wo�r�,A�)��	�-�Ε���oj�H4�ͣy� =�	cv�	{S�(��B��[�kz�x�h7�8nAЦ��_�A����x����EI	�`N���yW�p�=��x�,�`��K�1�&�����U>���C���5�`��$�ޫ�]J��W{6�i�_�Ѓ���Kl�H�V�Ga�u��7��x̱\���x1�d��J��J���8�z7yԫ&\<��@���b�x$Eue)����9���+����gq&�A|�4�\Z��*7�n2y@��f�!�1����-�/�߫��~�.0�Y\DK]����z���bm��$d����7�<����g��{���|�0��+99�R�Ҽv�{n�F��&�{b���[����^�}[ѝW�I�m�s�P�\*%����?Cq�1��	�����R���s��	�w�5���*� ���Ul��@�<��"/ω$:b#�-����*�X/�>�{8<�rؿ�	�]7�ņ�G�>�⩍/��Z�.����L���\d ��������T�]��@[=H�m��Fa�i���mfN��VA��v��Ҥ��s�dwg��!E�,���w"��2՗N;\hw���͠��.����si�� �3�������0��6#{�>�BJ��U5#�Jo+QP�h36�Sݒ�ѷ�լU�gP\�AmL^p�5�=��,�~s�<8Cx���e��mf+�3�`=�o+��A_˛2��S�:�5R��)y�gx��x7Ƚ���G;'01�n��mqN���L�-�� ^�e�E0	��(~"G6�?�T7��c\3/�����w-�!I�����g�-���t�a0Z�#b�4(o���O��>�7�g�k�3T��1K�b�_~��n�p�R֛Cic�$���F�hI@��r e�������X���b���G�[H�����vْ'�u��`�
. ��i����2`sL)fC�
騫?u?����[P�ˌ-��?�3ݜ�dl�W�1�0h��9S�%0s$��-�?~�3���SwV� f��ȹ�6W+�J��;2CgO��>z)f3��O���,dp�~7���!T��z�ǣu�sa��ZQ�xn"�-�z�f������T:ӹ#�a5j���>�
3{�n~d�[�����HR�R0�m��u�U�&�'fVQ�vR�$�de ��2TX����`X�	��8������!���z�b�+�hv	Ct�_�$�p��'>�	iJF0�%��ԇ~�Y�^��Y:�<W�\�k5�����Fw����R>�����%4��@OR~�OuuP�3ε���F+(�`�^��:Hh��c#LMe�{<�c�X!/ WJ�G�ɑ�wr�6������m�X���3,�v�S`f�0YR��v���s�&o ��Q�ۛ=I�'�r�E=w���������	>!C�f��� 8ZVȍX�]z<��e�Fk�a�|�� aΙԕ��l ���ڛ���0To=Ty��4��-?�'�h������\ߵ7�uspw�Z��6�a�
�W��9��e_�6o1�7���z��\�
1�6���֏!ڸʹ	:,)Wn���͟#ԩ�U1�}� z���A?��W�^��Bªv��c��ZZT[V�TlJ��s:�7Q��;Z�T`���X�����ҧ�:^��*�Ԯ���⑬=�Z񃾄ז�/.�Ｖ�@���%��Dg �`��G{n>�\Z��
׈��$R_å��.f5H_�0����D�n��1u�e0���N`3��~�u��QO	�k���MA�\���G��:�[�C�,��V��(��JN��%*�a�*�@Ω�����tI��18�1����.K������c�y��6�R���0���a<�
0�H�)�[���8�����u/\�蒋̚�j`���Y�F$5�#�k&
K��wn��a-�����At�k�a��t��m����|�����8+���|niTKF��K�+HV>���E�k�� 28]�,ʅ�٤��V�����F��y��qT�5���܈�r3�XA��0cR ���@��k^�~o�;�z����c�i1��4#n�B�Ͻ/�hēh�<�S6$Y���5��[nϡm�Y��s�C��Uw�q���m�g�;�8j�����ቼ�b�p�t3X|J�b�J�����hW�K���Ny�c�{�$nI���3N�����*[���6NGi"��(��aٌ�EG���ڴ��o�)��i��FC/�n�}�SRK�7A[����d%��	�0D�C{���Ik.��t28u�P���\P�]�
V�����,8U?;@�[��Zm�,mE�S��I���cK��h��7h��-W�ڛT)���6Y���Z]��l^���4�(7R��)ж?M��H˧�������3i��@�T�Y�jެ�9���T�#��N����r�Ǎ��TwLh���Tr+\���W�9�G(��&ie����%��#���"��q�X�I2(��C���\t�B� ���p������e}�%��@�+�&�5a��{�d��KL��ɣ�[_4�H4�C�A���|c��+����rWX�k8�tٶ�rzg�V�1w���Ӎ���?����i��=��Mj��@8�8�,W�� ����B����q^|!ݏ�'�(0 ��ҳ{��G?��w�KPJ��͞:�U��mv7ِ�J�2����qW;��p�I���Aı��N��Q|��r�5��j��G���t�����8H�Y�m���ك��`:s6(L�.GK�X�����:�۾��<͏�>��8�C�pO�bAjh��Q� L��eğ�]�!:)��:1�WX*7w7wn�Vt��y�bc�tV�+dk�b�w�ya��[�t��VV�_�/����OP1@�N�⯲��J�k�Q��B�M�Eޔ1���w���x<ؘ�!��7�8�N&e,�y}L���2X���]1f|���#�b7����Z\�5��Ű/��q�/��*��m�3�1ϣ��������m�����F�H��6��_0�����Q)��9�����lF�uT�	(,�	�o��+�8��g�\䖊:�����h{��g�S��/a��JLm�zzR"ƚe �����ɹ�{�;q�&gA&���<��؅�gX�n���W�S,���w��;X/�> /3,��+�CT227[
����[�H�VŗP�N�������6�B�h{W��+M5E�k]?kp9Ԗ�t�)�.Ӝ�w�`��V�) �띻k��o���=���<:�+��z���Ɔ.$��L�^���wH�X��p�Ci�u�?�J=�S�/c M��XZ�2�A���E�3Rw� q(Ki��8�5�,�u/�_�p�����u��ޯZ[��"i�'R^EZ�J��h{`�.%?�����#:cì	i��q��Fi˃�:d�$���OY�˱���@c��M�K�[_?��aՏ��=�F��f@F~(��P���#e��D������n���)��FH�{��O��˟��s���h⓷��"�.7��-�q�M������t�5J!8}��>�j�6]��1��aaC*�����Y�a
�7ûJ5��XqAg=�Ϋ����I���^|��|Ȃ
x%�Q�,
�(��n���t新��D���Q2��eKX<q� �}��g[��Ne�c���hλDh$&}LdO�)\�ޯI��x����kB��6�N�e��f��b����>��܋-���y