XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����d��O�r8e�ӓm�	U"�d�+L\�˳5�狻l�m��Mukr��<��c�����ǯ�d^���g�S�?��_2���Xn�%�*�5&^N�O��7��ǢV��6 ���f
�7��V���G��e�����BV9����_�SX��qyUӻ�\�ߋI����DZ	��b!.V���<�Ƀ _+��(	��EA�J�������W2Մ�'�!�9�p��#SR�$��	�A
�C�[��R�f��&-G�7��H�4��ooA���T׏� ��x1x� 	 ���t	�D�hIʫ?UT�p(%�<��Y!�J�{��j�\���6��z�׳3�!��+�la�>�����t�=��2�@u��mAh��ŏ��ݲ�7*����^���}�s��/��O�jM�����`S�G:��CA�F2�E8��˶l�"�L���[��1�%��
�l#Ϻ
���v�[<�{�)E��c.�]t�au �Oү���v��w�΁-��O�bL�����؁�I�Ws �"���5�.9=.�Iq@(�#� o��F�Gų*�p5Vy��.�#�Z��K�m��m�.~�1� 8qh���#���H�����_�5.z�!+V]Q7��g��=k5M��|W�K�bq�&??w��Fn����S��X�Yy�'ѝ�e����=���,�,v/�B�U�]G�R��Tv��sh���wr2���	-<���m�I�3�c���2���O_u�w-�Q�]\�" ���b�XlxVHYEB     850     2d0����Z��b��fU`��5�0�;�j���'��/8a_�@X�yz�m�fЍk/n��)c�U�Q�Ep�P�ݹУ;�(W?B�G�@�:�Ǚ��ӯ)��O�
ˮS���	Vp���"�+�[��J�2ܖOE���!�:�:)�A!<P�z|�h ��b^W����2�p��qc�`Uv
�����8�B�����c�i�q���"T�-g���)O�k����2`<��C3�+�q��(%��F��4Ƀp}�;E�ii.\S!k�P��	à�`��o��?�r�8�� 	H�M��ԑ��P��������cp�!�	c��VY^:u�+�G��D������:Hi
��,��O��5>�5����yy3�������Щ��t�<V��är'�Z\2��X�	5���Θ�RM)B2�C֮�}>"��Al�Э�'��ح��˞�5>%PxY�p.`�=ڗ'����a	���
~dg����$'�����!X��f�[�n����z�e{h�����_n��o`�X]]�����3=q�8F�w?�<��%,k,vU����5�@�J@��$M� �]ј���}���4N��}���!|�&����
�Gp��D�¹���P����I}���j�N�O��&��7�N��+Gi�?�~�Pϔ�l��?,NL�}�8�TM`���Eh�!mYv�ii�E9��������