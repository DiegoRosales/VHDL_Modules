XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���L��U�c�˦�ܵ�[E�uJ�t`<2��Hv<��5�������#ޱ-��|!�ܷ�n����[��]�08f$��¸��5��������c����J��v$�9���+��K)a*t�H��S����vA�\�_9bI0��`�@��u����'�N��v����D-t��fZ\v�/Z+5�)�h����-��K�jH�9��2�'�-Ca�;G�¾�p1Z�`(�3M
���aj�v��%��X}�k��M���i�h3�k h�ɨ2���@��=�+�� �!0�3jHT��v�P1V�[3��kd�A���E���:�4+P�\7��[��v�c�yT�1K���>��\Tt�!L���q���,�A�-fX��+k�l6��:�:�T����Qy]eiO.D�~�d�ۿ�(��\D���rw�����E˭"n�!t	���ԧ>���@P���lpt��(��[��e�5O�w��2m@{gb�Dh���k.7�g�C��1¤�h��b�o⥏GE�m��o�X�2Ky땏=F�5}������jp�����F�ě��e�^j^�{w��������
�l5�Z����Y"���a���R$m��B/�r��-iL�>�s�[�<�=�_���C{\�]�ٴ�r��7���qj�L*WJ�e���\���'G��va��<�H���e���>x`"(�_=��ن����8�Up{�x	�W�����m�"m��):Ԇ���"c^��V�	��n���.��E��{�葐��VXlxVHYEB    fa00    1730����� ��cm��9���a���qM[!�*V��.�X�N����v��F�M�����\u �@l�P��,G!�YwP<b�ҡ��e�6_�X��&ޒ3C�}t�<�5���^��5��!��0��l��᫄�����J����^70/:� uv"�t������y�+�p0@Z��.=6u�c�y�$��7 ����o���#��8p�AJ��g�gC�s���yHc�"�e3��c�2�=��U�&9Bh9��k[�1��d���!��/�O?yDT����{�h-8"/v$��vwN��|g ����U��	,Q�d��CC]�WK� 2��ފ�[���~�'�iBi�DB��dA��O/O�����6(WA�����̳r�PM�k�9�1�d)n�f�_[�������^ P^������o��� �{��<���i3�O�ZDee�2�r���(ȅ��1��2�@�5�W��s׾y��Nli����h�����2?�x��~���V80�#�r y �go4~���{�0suՁ��a��a������!BB��?���1���ˢ���Q�!qB�T�I��=�$�?5���Ӕ�R���E`0�OC��٦��A%��7,8i�@��T]�}�Q����Wׇ�IEs~���i�TM�o~ξq�)H��Š�I6�T�-����y��^��XJʶ��z�g�\�{�(򢽁@�q�������n���ZӮg�@���L�>�Qd����_��/Vҫ�Z��r������p+���J�v|e%�~����6�$Z���'��.ޙ���)2fg�حn���tb��1u�<���]P��_:��o� :��G��O��7M����sw7K\pwX��aȒ�g��?��{�<-j���iY	�����&;I$!P�$X�6�#׵���n� 
f��e��k.�h����� �EzMm�j2�c�T�оq`�����U[^�&#��+�S��O�gW�|R9`Pi�Wé�!���J�&C	���y��ҍ�����sf�HK�҅%:be�c��Yo�1� C��E���S����/��,9e�4]9<8�J����\7pt�"'��3��יx���{����� _$�z����vn۝�^{�$N��/W8_�@zƐyz@��U���|�QE�)�����]�IUGh܊}�%���C*�?X����T�F���N ��B��� ���щES�ETo#�2:9C'��DM��
"-��z.%�����լ��⭼vi���p�����,|?ŵ�M\D���?$�n(:������f�z�'=y�T�l�"yO���� ��5T��v���j4x3^��Σ���p�e���v����R>�����`����⍺n��[�|6P4��<�W�n�TK�^������[���+�!s�4$g��g�f��IW����Â��b!�)J�V�=f|�x���[��T+�P�C�'+0Q������>���?u�<�I\w}�h�h�/�k�2�G� ½}�KX~(zZ���1��Qp��k�V��)��Q��޶X��N�t�ͨ`K�Ep�!�_ )�]|� �'��)BJ�)y��/�uq,��(72�}GM�����j�	�*
�P*��������S�x6�7gӹ1(���l��*��,=�ök����9�eC���V��:�iY[�0�5�����&�GZcm=,�-���F���~��=~�:����쪣�'f �R$���3u���ZC��a�KS^�Q�h�E���y�:&$F!��5�)�[`�2���+�{�(�3v�$���N���tW��n��ߎNz�t�V>je�Bm��$cB�*t͐e�,>�?L�huqbַ���([���9s��3� b�@��������v��>jjy��� <Ȑ�:h�%ɺ-(se�y���0��-�41Tܿ���	�X�|��
���r����(�v��Q9�r�x��G61$�c	�L�_�ǘ:���ky��R;�{����a�t���ު��D�o�y��fw4k���� ��Ծ#Rd�3Ό�w[n���fx"��`:��#�c�G5k�����5��*_���F4W����Rݿ/�^�I�����a���ۨ�J �+D
�H�k�� VA%�0�P�Z�%�����i�(u�y��"`����s�B����TB��w�,e��ul����H>�����yY�2�98�L�����]��^0���}n8����ѣ�b��_'��\;��<��[�xli�@��Lw3m�6���0��g��V4��Z��{����K���P��E��'l|7*��/Vƣ�≋kV�'\�+ؽխ-��CqH��� @�н "|M�'�.0����E|K��C���[`|i�_�~5�$��,�b(�H��P�6��9�8��`ۇ�;C`�Sۗ����P��T���l$�F	�$�M�D�O���x��_������f+PݨRF{�����8M��y�t6�]�\�C�2�
co�I�:xy4��o���@�\s2ϟq��J��cy��&H�0�C�BE�K�;h��&PJ�Ɇ�w�p������;�.��5��M�lJ� �i�5����Ci~Y?z$���}=�F�ސ}$>����鋗gW����'��_z���n���>O7tX-Z.�;Q��ybI�Q������:��E�i<LݏB�J`�dYs�y�qoP�����4�1֐��P��ܩ��H�<��S�"#�@�~1GA1B�1�+PiQ��nb���.X��ƭ�Ye�{M��İ��zW0�
�y`�/�/���{�� L^.�6F��B�J~�ɷ���;l���є?��7ى��M& ٞ�e���|ZL��q)��^��m�]��O�v6M���R�/�}�Ecv�7��ez��܇��<�����g����!�J�FqS)�ص�덊�&V_�ԅ�q��:�
ݙ����B���Y�9�z�δ�P������ۻ�z�s�P�*�;�g��Z�BH 9=zR9�U�m`��1d}4�%C�WP�~�x� �E]��Pb����X���,X��2V����cNU��q��C���_��ˊ�=�]+8Ӈ Fͳ���� T53/�g$��b���w���a�2�~���#�c={=O?�V�9���H$���>���U5m]��K�w��Y�/ =��J��һ��$�ݺd�6�*0Z�2@]C'� �ɉ%�˼�P4u�a��ͩ��:,�/�(��q\q�}>���O:*F�
�9uS���2x�r�9�D���-�6ف�{B7,=ƨ��D;Tݮpc����=2��`�޻�:�U��rZ��mk��}=�3�\��x���dX�&���]��}0��hW`���Q,�i���;�T�
���-������"�_����%	I
�V�)��� :�{��&���KA�XB �$_`0�[�ɂ���oV]"�9��KoT)�������%y��(��)�n�W�2��\,ry�AA%Uū�)�X�"���x5�to(�f�/y�B�=��|jG��j���O�v]��ϡ����˘�8���j��x����n"����o�Π:�1����Q��*��>P,�=qX*����@Ӗ7���V�\b�lI��?'1=\�l�4v))�ȏ�\��'k+���>����Us"��p;=��ܚ�9GŶP_�Z	�*�#]�� �$��{v[��k@~�9��5�>�j�u.���Q��'D���c���J�W��[_o��lZd ��egD�s�,s8����T�&1�
J�o�C��Zdn���9sY�Q�ĺB��*�ͯ8w�t��?q����?/#��ۺ�%�����WmLL�!a<��tr,�/�.�،��i9�bO��6�m^?&�c>*.�/�9� �(�����,�/v��y9)����./�P����I�|y��E3ʫ�l'�����b���8K�U����^e"��|��N��MۺEo#��u�?	&r���nq��evUJ�Z��?�i��h˱����.x+)����k��f�߷�����nbՕ��EK���bi5<[�b�]���Z�����O�
��H�(W��_�'�,I��(}��z"��G��G}��[9U�K-="�}�1��I8⡚I��%7���YL_�l����$^����FyE�B^�ò�%��9I�r�������H���-�!�o�W���Kr�|W�3<xh�=�xc��/�Q�Y�� O�[~����5ڋh����\&��"�pG"��rx�vɩѢ�x��D�T��p=3���#��#yLA�r�[������{�;��ګ�U�y�A����\ґ��b��hB5�l6�Y^R,'m��O�2S<�5?�8s���4��sd�9K��5���Չ9O����tN�ɾ��1�1 G�I���#�~����Sf�6T
%���W�~L,�(���)z�J�,x��Yp#�ס�b��)��5��Qc��~�3[�pжn:f�~� k��Q�G�u����%$���-=<f�g�z��as���K�waeE���#ףD����Z�\r&E�	j�cX��@N^�Ac�ڔ��|Db��^f���Xe��._`���OQ־��o�1I��g�/5l�l��"�����_.�O@XG�m8 ��`�ہ^jPƨ��1Pa�#I*u����`���_�C��R��a�r;ϥU�'��$�(:�Mi�������<P���0^�Vʄ�3���;ħ �r�Pb�߳���o$���<�w0~/�C��	uQH���ߥ�*��*
t��c`� ��<�I�k��g�v�㊠��B>WM9�,(6"|�|t�I!6$y\C���xx$6ҵ�t�Ό��7�8��*W=�u���pu#����m�zH�l�,�����F��_�[Ou���L��"l�?�7�5J'M5�[���3,��aX
G�����9���euv媉qڐ�����|���~a�߮;fy�������o�T��1�?Qrg�_������#ں�D�웱%�5t͙Y�P���8�9BT���NM�d� e�+��.�
� �Z+��e��q?�c�Q����"�cx���j�$�� �}�@H�0�g��Zng�����B
��x�_-�I�@�CY!�}�He]<C�r��M��δ@̚���4I��;�?"j���&LV�[Mo�֎�D#o4 �L�j��\kw����6��e#�~u"��82o��wb����s�]�$�C巾B�yC����o��+C�����"�3��*q���MXY,���0`�ט?'�d���%���G�W��R��ʭ�z����歐��.�^�Y :���'�)e�e����t����U{sC���
�9��X��tj֋g�A�;�ƑU˴7�8�?p٬�)��Msy�������~Ο/�L=*�>����Z@e�I2[�l���Q���Q�[������ t�ӡ�����R�M̒! M����BY�[�;�&�iR�OK"A�k����d��f��|�b��
C��ʴ�;M��GbXK�8��Uo0\�5Vk6�'��j��,����E%���-J7��v�y��%��4
S?�W�����r�>A�.yV�Zxda��N���u!�H=��Ж��6���H�	r��p�=�Ns��eT�7?.�ָ$׍��*�B���Ss�$Y����8y�����N�K���$V��<�?���l^��Lx��=�ܼ�)R�f��*�W�m�#���B�̩�y�˒��RD�c��%�Mq��.j�f7�2�� �K����
�2
�R����@� ��nI�qy�DQxUխ��[+[.��8�ϴ�0~�[�)W���1c��y�P�@�G.�i�a��_XlxVHYEB    fa00    1d70�t�B�@3<-�@x�I��A|��eQ���b�ɳܠHF�A0�m���F�� ��v{h���G���/�3��k���<-����j�����$e���C/1�����$d��~��jdP����S��ԏĵk���~��ǅ'���
*���*��0.��������|I��d��K��=��~�WTs�9[��rg�*��%#�Ӑl�M�\��(Q�0�_`�j.ֲL��lf\K7�_�̋����П����,�c��a8:R:��MCK�0��R}R\g�V��S�F�]����7��K=y0��8�0sP���94O�l7 �ɼ�h��C�(x�9#9fcF@�DՀ�y�e�' �z1�"C-O���Rr4�����!�^��٤���w�]�aL� gn�a;[Y?�����H�r!��u.P�ګ4�I��R��z�!L/F4�I�6A~�Dɶ����-�nt�t4�i��*��i�{���X�o�Ҋ�WV�0 ��>}��B�*w�ƴ���V����y����WI��<�J\�_��
^��C�CR�`���=��� V@�m��y���N�t�����{�4���虵n^�V�9^�iV�(Q���yg�W��嚻 c KP��Љ$��(I���ZS���/d[���l!�PKۡm�2"]s��n���������jqB_Q[�|"~�U�o�cM�c-C�p l|�/�Cq{�%�ڽt�Վ/;sz~�,x�Q�b'PD\"o��K���,
�d{~�2�Ŵ��&�'7��T�2�^���vi�i����|Z��[�u�
�$��M������YT=�!�1��)˦2>J�qS/�i,�8�z���eQ<�Z���-�è��ҥ�D�D�Ζuuڒ}�����u�eN~�0=���j|3(ă����Y��\�l�ܓ
�J���s�����g'p�s�Q>��6��u��XgU�Y�z����b��`O�%��J�|$�]1"E1��:X��/H�ڴ�C؁�;_1�c�ym;���qX�N4���Z�4����12Px�56�A��5��#f$}��fY����K���Ŷ�����8�a���H�3���&t�>�X��1c�׎����d
���j|����X����J1��n���,�5��n��%�,]%�p��Զ�{�S�'�R�nJI%$�Gkg�J��R��	�0Sh�g4��8�h���z�L���]��/oo��i���Q[��y�1������L�=�%Ӊ��_A����)t��U�u���s]?}�*��uf�,\�C��3���U�����sC£�Tߵ��Hg�!V���������b��\�X!qH��	�`�(6H,<�tq�'��1�P��Z��[:���0J����PN�]MfV��q�[F���k_y)H/��ݧ�U�I|�7%�m�{�
e�>��^��ׄ2����P�G�v0Z�Х��uPW�_���C��G��LɏLkbl �p�Y�z����R�(~�ű��E�բĐC��`mV�J8�Z�m�Z���3O��x�@�+V~�T���>�BPO޳ˮ71Ǭݦ��ڔwP�Ppf�}��4K{�e��
9j@F���V�dH5V�9���L=woc��qX�NΔ;Cp����GmX�+����S�IN�	�W���4�-��'��vDܽF*�U�1��[8�s��1JS�yS�J����Ҽ�`�]N�p�t���֯�{����=���P��<ެH�����Yn��6�dԽ��}Ub��K�$��\���,Uj���~V`���,Aw��d�����@�u!���4_�P
�q�"s.�'�7�9Ư���g�*��]���0�}g����^�
�&����q�j�Q�6��B�6["\``v�����<ĺ	2̌��+����ڴd��b�$�,��g�EE�m'YY�ӈ����m�ŤJr���/�j���������6\�`�:���A!��;Wŗ�o�jK��5�	��և�����չO����`�+�V
R���2����k�d�Ċ�|�%hUZ��rTp�C	5b�?g��g���,�Q����Q�-_Oj��L*���TV}�'���_�|�����C���/�[�q2>bv�R&��Gh7��d��2�-d�Ņ�U�h ������o�" �I�؃�E�[7H���Sd�bl�.�(fᣜ�dCwBYx��Z��j]�x^��
�+�0��z_���5u��ј�� ���~4>ωv��^6<�+u�Y�!]
��95�C�k/lCE��?�rQ��X\Gu��P!���H�����J��T=]��
	"҅u����!�8��D�����)UQ<��>j������h��ǰ��`��v�lM��.����{�^Vq!�J�U�6߅�w�%XJZ���]�x�x6��þu[�>���D`d��|���ٝfst!���h  ��m��3~n��?uLw���B��s���]9#qɆf��m�Tݴ�� S�Q�P̶	�O@����<�|�ux� %0C񫸽�F�g��C)��r�`�� �gd�u䀲BP)hHⴏQݣ�q/��<[QP<U?��nc�2�"R�2���t,'�����K#N�5�j���r���l�w�n�����xt�O����=qz��?c����J%71 ����1����-K��wu�W���%s��#�|ـ	�����t�L-����Ĺ�?8D���Ւ�e m���ڒ�5"+�%��%S@��ԠL�
5�Ԇ�GM�-mĚ���N������a2z�E����p+��&�ǻ3�w���_�*�KIX��]���
�>����������ü_-v��´TC�d����Eu�|d�k�+p5��$k��J \���LG��`���& B�>rg�(rL.�s�@G֠xO �t�0��P���#��|j?�"U����6�~�Ҭ�C�)$ej��~0bF�.Cc�R��|X}�e�V���B#L�Xg��e*����|���=_��d�#c����;@�-�n�W�zx��1Ks�́&@'�q��r|b��k�4�����W�!X�eEM4q`t����v���������wl��z���6͖���M3�9_�Ie2�l�A�F$_�������%��q��(��+}���RZ�]2G��L-jB�&�(�L} <2A,�wE�m���r��6�y��3b;��^�\�Զ4T��bi�Apŷ;�fM��?���p�#���W��)�Ю� �.������"J}jx�Ƈj�2@����{� �2������k��|Y��ˎ�d%<�P�`
{!�<���#@��|k�ĵ�͗���T-��%�'N����vh�
s��̕e��Th��m��|&t�-;Df_�#��r�)T������Ý�~�Ն��̻d�5�C��;�<�nWȓ~�!u �e�ǆB��f���m�۞9wn��q0H�X����ǐ'���Ӵ[�����{�x �qĐ����Ƶ�=;A8���G���J��ؘ4�㶃L������N{�C97T��b"�K�Wٽ�xo��O�}�o 3�ԁ��X�ll1B��<lJ�Q�;R�ΦIEá��Cm[�e"�ʌ��M��,`�m!)�!Ϩ�R�A(0_����B@�R|�Hɇ� ^ 7>%�2��/���]dc8cK!?��n4�7�#T��E�?�~2��cZ\�&t�jfCuۻ�7`����d1��4W��~1Cd���j�-Ҁb����E3���bL���`V��H\(���2��9M�0h3�\��p���O��0&�/)�g�K�ӂ�U�V�K@i���@)�Je�2��"�q"������������ ��Л�󐸅qHO�IXrE��)W��p�Ґ)�<�.4�f �ӡ��Nj��io7�ᮧ�"�a���K �h����4�*�J��
�����D�&��������)�>
��:����
�#�����B1��M�,lV�m���M�a�M8��SJ��2����:��+ �:3��7/����%/��/G�!��oL���u��jKD�JU\^�Y�D�Yހ\������XQ-뛬�	xE#E����!��	-�lbX�d��Y�h���D�� ~�x;j#I"$+��I�� �1�MC�@���u�m���'�z���V9O*5m@���QI�P��j�3�G�¨GDEi�r��v�{e�n&)�'��#��h�c��o�n��9O)��$�0"�٘���t"r��.�{�sG�HC�^��;k��7�q?����c�6�I��w�`E��h~��ʨ9:UE���}�i9=؋
9��N�����b��ҋ���|�#�����s;�S0�9�~������f`Z��'��Ir�u�3󎾠fc� �TP��سN�#j�W�̇U�՚\~�N{z������\6�)J�y1j$ϛ��ļ��v��w�_����`�ڥ�����I�Ud(ǉ�k��$�sG3>�<����z���:
�0���6�ɬ��tV+0(�ɞ��O�V���>-	y���2��T�4$�&pAd�>X�o���isK�ˠ��aWB�"�_)J�&;��i�p�"NV&�W�si���@�DV�\!����C<$ϥ41�����4�q�Y�F.�w�;�KN=�"����Q@���#e�FH��g��Cn���*�s�l^^i������>O"��$����$�$��u���>j<S���0���h^}�k,WGiN>A?cpݴ�Ҁ��m/$s^�kLЕ�C��#q�\^ڪ[��<4tHa�V�ߋ���J�@��uP
j1�{{T�.ɞ�fT��]5,��D�@)��\�YL󨌐��q���Q��n�Q�xEHJ{xI��2�~�De�X�q5�gU�<��wS��{G@�_#���E��|}]	E��v����6�b@� S�S�I#�f����eQ������Wu)b��?�^�쉱�B�ƽ��z�����Y�D����  h:R/^�v����Ps���y���Y����-���j|R�uJ�v�M`;,����

H1C�gH#גi���(�]�¦5_�0���Ն�ya�J���
�H�e��{>MjHZ!�HR�4��&n{����6D+���_�E'�A}���� ���ws�G�*|������>?rX�Vc�����5���+&�j��US���4f��R��AZ�f���;��x-���,��ix݁X��izYN��-2��W��H�!�U�'��'�I�lԿ�����4l��}�[EN�r�Jo-os�w�r���kEf���������/,�1~f�S`���DJ�)��[@
�:"û'�?f���A)�B(�`��/*ŵ>��sןA����a�Z7�� �X��4,����.�!�	�m���|3}�rO<L%[���r86���/
�)��a���0��qwb"ޔ��H<U��uį�#1f�v�>�E�7
Sc{�Q�b��-'�߫��<���B|�#��]##�g)N��:�����:��c
5�����0�b%TfZ)���-c[�!�iq{���G�1�qө��Ax�$��N&��P�L��	L����FF���.>��L�&���e���_42�2Wn-eV��e� *��7�CU�ˠsF���3v�x���Qt��	�^y��==���f��!K"Q��H.�L�vB�����մ�� {�O��:�!
_�˃_�CJER�ަ��t"������%t�*�� ]�CzdE��B<FBd7XJ�/�ӝ�T7��\g��׮��J��)�Y�g��˞;�t~���>�@l��	k-��%z�Wۀ���Nbb�p.�5	(Jq���o�S�@��J�s�*�ؙ�cںr,n��j>f�Ktj�҅�~vi���FIƭ�m��y��61�D�� �
7��VHj�h�p`�,�^"��2,Vτ�ľzq�A����+��?��()������e�|��C����x��ѹG�7��?�.�VH���T�ӶC�B��c�>�WS~T���}k�w�ȆM��̎Ċ��M���8�I���,�^�r��7����W�2�^�G�|ђZ�əLg��s�ZTu�;εǁ��f-W|U�ҭ�N��2�XK����@�M��nO6�q��;��w�4HK3<���D��Η��`E"��Hf�
=�x�q���鵢�t�O��3Te�2����f]pi�18��Tk��\"�X+�����.�iS���v@�7�T�h��\�M����l�Y�vb��[BըMRt*?˫�B�a��5Ih\�ass��9Ҙ.����D�H����[F*��X%��FO�ÿ�91���7,F�0�Y�m+�'��v1�:ʎ݊�]�}wc.����K��g�N0�b�����&�Y;�O�G�AD{�k6X�YOe�E��+yˈ"2�M˒�N�X� �/��krڔz��G⯃"�f�L]Y7!�\��4�)ٜ\�j�ݯd��N�8RE�E1Id��v:�aC4Ѻ����i�$4�L���@�?��0�m}�*�5��pR+N�؆׌��2er�zc��@���%�=ߚS�ut�?>�NQ�#�����
j>:�H����qW�--�L�2�\S弋b�|�-��Q�� _4p�C�q0oJ��w��x�b�����JC�,������ãS���]��t:`�&�RGZ�=�c�U�*�H�u�{���U�5`��X-��B�o ��v��h� ��D��[b���2f��u4���7fANQw�l�GW��
 �8�T*��U.ˢh�:w-u���|�Ah���W*�v��Yy�kX������f�V��/��u�di��xqj~�O�BLY�֥�� >�SF�+�����yY�������p������I�G�ι��wsw���7��녧ϐ����	p:��~�|���W�e��&��nVu�5�{�M�ˤ���4���.Ò��8�! 71�_4Q/!1�w�1���_�9
�_y��#/n��3��o�R�Z�z�DͅV�9=F��� 1����K�r��g�7���EH\�0�Ԩ.b��`������Ø�
`�T��jW.׊�fZn�ӍB�F�^���E#��"���U��e���4mT~�s?��. z�P�#�|[��b��r��gl�'"��6���z`I���k°����n\�2jK%a�s� #��ߥ�O���"�i��WwC�DɌl�5�?�"�gy��Cޮ�KiW"���lVvs>��^;?9#	7ݾ�ۍ)�������t-h���y@��t��7�H'��G]��O>I}��c��f�Xe0�i������8�5ݣ�$�	:5�'�RRuB@e����N¸4.�`�K�z���~a�M_�������s������a # �E%��@Yӈu�<��w2��������C��%(��1��p�3���E�H ;��I�^�~Y����;���_�XlxVHYEB    719b    11f0�z����V�z�%E@{C#z ��e7�ɗ���l��!#5������w�`k�v��
��̳_�a�@C6)R�!#����8P�H�>�kY����|���eK��)L�q�>k���8T����	���r��D����~�"I_���o�x2|�~�'�Ɛ�L�|+	g�(��[� q
�� �doҍ=���MFt�#�AP���v#D���y�1�ZB���X�'�P�Y�֭�����
;����I5�pϖ7@B����=li��҉���k�N�Z^�Ǒ�+�s7�C���s�&Y.��9�=}C>��0^���y��L�~t�ciۂu�khkj&p	:'*;2����8��$����u��"���w�Žm �*_��m%������"���3�R��L(Ʌ�@L
xN�j\+p�-S]�Q<i��7yi�^�tP$��i��e���9��;�u��(���g��n�yn�[ڜ���2�bJ�U�h@���aC?�V� �����B�� ���+Y%��mL_R0�W;XD����A+or���p���;��q��o9)���\�D�I���C� ���F�ϔ ys����K'쳣��i��ʕ����$%I"�C��M�3T�ܾ�2��+�6�E�,�58�$H�FWWOZ�����l��V�3��@t�?�A�?�o]Y}*S_�ٻJ6^��_�a�+��|�Ҷ; ���a���p29��2~C^s�L� �?e�Ζ���xq����Dhr�U0E�J6��&��9/�LD�ᫌz�z��p�i�8�V�No��:Ѕ�-��-g9���+y��#)	\�d�Jbn���|N�oA�i1uJ��KMd������iA�,���\CB�}�dڲӀ���P�	�^I�w3����/������&�����'mF6ǬB���r���J�ڐ�����*,�^��쥇|w�v��G�,C���5��c�	�*���5�&A��m�rU�ϯ�G�M���>�]�N�ڇYk5}M���[_U𘨟� �1:��`��q�	Q`k����=�܇�XDa	s�T5�w�\A���Ɔ,k_���+�W߭nN�g�47�p�d
�*`�j�+�
�p�*~�X�c��تo�0)�����i��~E �S���C4#nF�;U�d�c}�j�yL�F�����#��vtO,kLA�5oo{�%6�kKT��Ȩᘒ��^&�4P�,�R�"�?���`�('
�O�컽Gv��g�vNy��-i��:V�C�Uk97zU��08�n��5��!��0X�P�Z�7�����v��;�ߙ��+���%�}���)��%w�Yũ�7�N�m��[���dLG�� �C��Š2�W��'^��(.A�ȍ^c(7������xԽ\�-�l.�L�����n�}���*�oR�A�g���T�����'|���j���׉��!#[�ko��-8��������0���]E���0"<�)�$�*F�o�ͨ��1F(T+�`i%���f��,��%/VW��bN��P܂�ͽ,{�P��~��Ld���� ��7-�����^���Tˬ^Y��x��|�W�h��uNEe��9�E¸��3*�2���H��������.O	�h�GD#�G"o�-�Z7�s��7�?ֿ˹;~�?a� �-�D����l}�:G��a�2u����q8�@5����7��]쏇)��go���1.�y:�K���7�eF�&N�,Gq�R�AG�ܐA�':(�Aa����}%$'�EPX8&�[{j<Տ^����IS�yUH�P�x�ԕS7�Ďt�h���9$9���U������ԳYo�&M��ں���Q����T�+����vF�K��4�H�󗄔# W�w��^���e|��?RKG!��Sy�9��&�9b��W�'v������k�]Ay��'�WA����l��K�WL�˭��1;*\��'�<p��m-{!�Xt'=�]����;c��+ ��H��%���?�>���޵;V��K�x�����<| ~�;������ ��x<H�t�
!,:h�p7�+5,y�����h���̚�t�o����;g8��hM�]j��ǡ�A6?�("���"ze�>�{�	Ք>Bk�w�^�+c�I�K�V�
w�z�Wk���X����}���#n�^�$�+[�S~�������;��H�t�:�U2	y�N��l=�F5w�-fRr�7�|�Ei�w�\�+0��Qa�������H�2�a?;�a�뼔b�t�/��y��~{�,�縕�F���C ����%�9Ζ��p�49Q�"i`Ӻ($��� �T�%E��t���e�@�6�����i��'<S��|�o}eB6�Ҵ<��c*�4��cJu
9����j"��d;:�~Ȧ�Y��meS�!'�"�s��fak��V_�r�b�[!���C�7�(̼Wq2��_.G�(s�f��gb��A���]�%�.��R��36�>���?�G�Vb��đ���O!�YOJˏ�vk���ɤ� �Fv�F5��śnt��?^���B���n�b��)he�)U���G��e��X(4��˜)��*���G����j%��HS��V��ი��*��i�a�u��*,_8�Ok9Ū�W�4����dѷI����iQ����X�3κ�,�v��� ΔY��V%���5'��u8�u�X�����/��&@n6y�ώ� pU_�Y%�,�UW^	 -^�D>/5�ѐ�5��T�=�te��+��[�W����؄~�P;�N�D��ޥ�5>^2�fd��"��ӱ`�k*�,p�d�dy���Ț��G\���q��x�F�ה�H8�S����8�T���r&��9����&��=��a�c2���{����r�V���
��-_���G�|�+2t�V���X|'�=�=ɚ>6ՎU��s��HTaUNu�����(� ��%�d�}��^NQQ�0IѬŰ���(����<������е1!7 ���-�֒��0�a�Sf!�Y,�<��h�VxϊE\�x���h5�c!G���!��%W�C���u��\2��G���N�ސ��\@5d�}�:�6Lm�h����0��>�&i���|�rG�r����yP�%����S],����h��+c25��Is�=u=~`�-K�4qօE�����PD/#�w '�߱��޷�ܥ�Mbc,��F{1L�� MÃ�<����!(�_2_m�#5S��� ���~S�� ��c��處��r�#*���+��|4Q3cƗQvVy)��|}pXx�$_dW����n���>_�[#��J�Z8؃��;�=�@K�� N��;��1���h�}�l��+���1X�3R�S ��
��٠�K��]�wٌ��q�����Q��ˡ}~�rEŷ�d�o��Spf�����1Z
{(Z�:n�)�뽳���^w�U���]d�U3��Bưfk�`�ee��M\w 5�n0�f{��qu�_B=�a�$'�#O	�w�ϙR�B� �Rք{J#&����"����&[m����afT�28362*��^���`�9�D�;�~�Ubn�e�O|;��l��F�t�w:kJ�&�J�yp�����I����c�����ʍ��7�;Wp8����s�#w�3F�ol���/@�+��,.P����6o^����͔i�������{.rˣv�f��3�@��5�x��YV�?�n/ߓ0q��-q���YQ)�g�ׅPg& �4C+�pTZ�`���Y����V[d+ǉsڦ́h{8�t%�}����V����z�;��H���.&&m=�C��gT��ka�
8	
_�(u���eo�&��աq�F�u<��+��"@e�P�$P�S�.R7�r�~�kM��o��z�u��M������O�D�.���{�FS��r)<��dόbm�K������nY,CGg�@A�i5	V텫&�i��G�j����o��H�g��6����9�.Xbuq���VS�{;��1Za�VT��) >ɘ���x�
�K��LZ��KKiЫe����#�D�v
C�(�~:��D����ͷ��9��I-��
d�ɦ=r�G \x��cj$45�ڡ�9��Dg���o�����&�Ʈ�j�����U�C3Z�o��Ȭ�{�_���r$�����`ځ4�fs宮�-amd5"w]t��RΰUq��\�*�S}�&��;t���[�Gg�[{퉔��l��e8�Y(E�#$�~�7<��:��uu�5	�o)*���1�G�9��vul�d6f���M��nF�@��/�����K�
HP��?ꦨ#�a{]k�F���WEt?q�E�TO�ε�Z޸X��I�vDm��'zs$G���#:��T���W���1��-}W�'������Fnj�O���A��^�[5|�YP}RZPӞ:Y3��\�^��2X����ey�5
��s" S�)�F��ą�DrŽ5Է��+�!�M��+�}+i