XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��	�v@�\	�^���XߡJJ�_i��'m��zsSf�]DJ �C�Y��	�VpL��[B2T~�i����&zcN�ji��Z�:��x�=��&�k��A�
lD��'�c.5�*jc[9�0w��1k�e\��f������Lf���<����\�Z-����L�D�RݒY]y
H
T�*�'��C���23j��|U���"��L��5|�9��uh�=4[�i��m�]6i�%p�N�>j��='�Zփ�U��ru��W18\��hUD��͈��aL�c��7�����Q��Z�N�c��m��-��w��F������,V��J�M�(4'���A �S�-iVW�0&����܆��dz=_dfVߟ��Uv��<�P
�� �gGL����O�Z�M�ю��}آ��х��7i�]!���.}�g����,��-a�g�F�hW:DQp�]5�dE�u�6�<����0�Fk-c��Q���4��UB<t�7�ydܚ�ux��KC�m�r�!��\e�5��f�֟�A�r/�[�-ύF^��(0������GZ��Y�Q���+�s���/�x�PS��I�3ڦfX.T�_(���w�����`�16�_�qޯV�#1
�,�a��E��� {}]=k| �{Ԡ��\@���i~�8nxԧw���{��*9�&>�ǒ����g�	f׌��$�B4\�f�p`M�&���6������.H��@A�!�\���ӜC������35��8�����`1?{��=ه�XlxVHYEB    fa00    2ff0��O��5�X�Qց�p>�@�\kN���Jg�@eA�ϮO��o��7]��n�t�HpwBuט���H��-��^<�<�Y��9��l'[�"Nm�%���K����s���'"�Jl����i-��&�F%�_�����C���}��� DoZj� ��I����=��Kn���x�BU��d'ǈ��PC�M�*��K	��%�p[�"l��FF���俸�sG�z]֨6MJt���&I�V#���+q!�dQA0�t���]�� ���6�=��B����H��&�ߣ���w=�8Hܘ��gЛڽ���p՜��������	aU{�{��Y��pȈ�q�C@:�mH�wzm'��WJ&G�����e<���A-�[s7{>&�����obfW�U-��y�Z�,��)Cet�CK��٘F���>W�g�, ���'�)�-�ky��k�J��	W�f�F]�UR��%_�%����	�F�47�����1;b�~�j�	���TvF�)���FB�����ִs�M�]��t�M1�kEǠ���q��L�.-7��
(,c����s�t��r�-Yj�s�.Zj�{��`�j��k��P�8\r�(�U^���6H��l�8���kà�,��x脿8��r�3�
�tI���7ў�}@V��Ӧ�M��y�=F%X�'6-V:��{�by�
N�y�P��s�Օ�*�0���+H�ǁ�{�j�P�4�e���A �~��B֢��H���n��4E��a6)F�c��ؿt|q�>~=�H4�(J���H�Z�i�um#��!s,�ݍ�M�Kx����|�a
�曽��>g����3���;�m�M�`���d�g��5�4����܍�̘k��-r�0�3����k[	��.#q������v����|����	�LE�h[�x����"�bS�������bD��-(t�篛u��fl��
� �p[��l�'w|ח�5�T���8n�:�k��%�i$S�+b!8����=�
W��ٜ�m�4�q��ꎸn�a�� �ɃX=-���\�c4��{>�Y�%��`t�#�(|�Pt�%� �F1�A���75QM��{*'�k7���a5�T+��u^(-&F3�m�:�$�e�Q�K�+v��r�8�0$��U�`)rX́&k�px�5|���4J�>��(���8l���?wK����Qp�{�R��p��C
f��V	�ǣ��0��y�mo�*.�1c��BJ�Ⲧ�����6��BZ�2;@�5i���Nr&z��wd
8�����?���fe����LF���6��.�,�o_,!ڂ�S��JG�J��h7����Qaʗ��^�Z�ޝK.:�$��p)5}�\K4y˺'�)Ec9�ίүWH��;S���-('�/�:U?3Nf"�n�z�q��аRCA��z[�Dw�GZ�+(kQ,�  �Y����8\�awn�m�)��y����L�	+凌���F�c�� 
�,ۢD�i�&І��Ĝn�m��9�2J��:������?��M5�wQ���U�Z�X�&�Q�=%ւ�j���E�ڣz�w@�v����� ��F�I�+R!I�!!U�+�+�j���GؚR�e�E3��i�3 /�+%!�&�����N&%}Ώ���� ̔f؝�8��a�֓����_�f�"K�eJ�/��r�R8�H7q�۬W|h���5��3��kV�Q5��qO�A-�̕%]f$Y}-p��v��C�Zriq =v�F���-��:���=���Oz&;<��/8����ZZ�iPi��j���G�t�YV�X{ $}�����b��t�G"�&�{}���7���۟�ٰKT	H��Jܵ41�z�:O�9J�Ԏx/�>�����8���>�T�t
mYS$,����_Yvl�@�+�08q��eE�%S���V��x+:�+*�a0�_���w'H�I��X��_C���U�����Y��g��^�z5qW��-�+��#%gmN�gjQä[5�xj_�y�U�*j�茮�+�,'\�샂?��[^l�k�e4�a>�ao����KБ^{V����:��a�ML*�S���d��X����lm��A�N�W���N��]�eو���.{�����)��~���r�y�ۊe	�9 T ���.eg��1�מ�[M/��!��n���7)��fL�J�gM}t��Z[�:>�ԟ�RH�������r�(��ԗ�r�2��o�o��Hv�ϡ�V�4�����'��i��AŘwds\ߋP���a�y]�6)n��[oz&��ɴ���vs\��E��>1�1��r%�7��tN@�d�$kU�J&��Ǘ@P����O:�L��WjE�:��P�j�7�������>O������hv�:Pj�F���RR��u���*4V�:���d[��{�o�L��*ͣ;�l$'�y��n,3$����!�R�>�d(o�.AX��[����خ�AggbB��v���y��Ԥ>/��+�@���7�520��[�8��%��#7E��:dn.�׋N�SsRĻ��q��r�얒����BQ��WU4(�c��uC�A|��Y�Z6��T�vtiB�4e��Cpf>��p7�o�q�В,����?�p[O9�Bq8�7� ���2�����;�2��t|��oR�����)�z~)]L�.�3�Z� �M�<E�fQ���螒@��0yH�S�%FI�?�@�aR��J�v��hP_G4�6�!oٺ,1Ly��
HWZJ^�T�4�/1�P��%ԆtShcD�}ܵD�MH��fĄ��v��Чv��X�ۥ�
���q�.�~l�/H(���I�5����+��h}L\�?j��(=�vj�j�ޱ��Z�Z��_�;��h���N�X��\���~���h���y�
t���!X6�dY],L���F�}�<�t�)o�$��qD��V,�G;�����*7�F �i>����+�o���ի��qo#8���i|+��7M�e����q�.'�һ����H�8����%�Nj�����jaa��f��[�U���!}��>\����G�(R�R���HwՋ�	��۽<	��e�c��ǉ��Gb�2����;�x�D����n����m�����L
��8�3�< '\eS�"�z��X �@�Y�*E�ǋ{�/��s�����us1k��Fb�9ֺ,yYR�!Q�447_���=�n^!��֑8~q��)��Cd���&�x-A(~2�"D%8�n���@Ot�%q��^�/ek��PW<�m"\�*�(�?���B��aN���Ȟ�y��W�!�:���7�]�eª���9�4dr���ې5��_�[N�����>�H'���Y��є�9��K7����7�om�u�s���

�6:�)Z�����������Aۍ�&s,�����戋Ϣ@�2���h�ω�VXVU��Y��e��reԂ!���!�	��%���v���Pb+��u~�����1�7Xoe	����9���9D?�)�<J��^B/�C�<b�O�ݮ9�T��f;��:����;˥{��ݾ�)�����"�y��j:��Ae����L�'D�-��v'|�Àty��v�E��������G��,3��(ą]�����P
�ܭu�(�=��fd�rGh�3��GnˊK�k�>&`b{� 5*�z���3�Z�4����J�D���Z���,�rަ|V�
����񧙞�.���@	w�m�o^�
O.c��2��䣈��C~����1��
w8�l�9����v<	Y]��4�˟��ŋ����wB����Ӛ��5�"&y������j���T���K�'D��[�H4Nb F����,,�{�{nK�9f�&-�;wZ��ЮbX��eE�z�o�����&��pk;/�����]}	�'{���_U5?�Ef��11E���D;�lf�V���ڿ
V)m�?x���.���4�%
����P㫸+�v��"�$2JA)՝��z�mJ���@�c�-!kM�~>1yͤ�t���V��Z�N��� :�v�@hA=�*���:Ű6Dӥ��ƝOlm��|����kO�M���<���n��a(���H9�&^*�|0���"\���z�Ya7N��Zs��v��5m@�Q��FR���le�X�9�#j�>��b��u6�)��
9�bF�6���J>��gB��^A���<�2(�����8��wO�>w�)l�:8�
�����ߕM��}����ʖ�h�^m���f�B{�����ô�爬�6�xp����w�I�qJ�ɺxI;0�:�x!3�%�yg�N�*۪�@����85�:�8�8M����4�Y��~���2O o�o'��'���ɸ~B�����;]~����T�\�ǘ�K�6��-��1�B�ꃔ]�<�����:�H�#Z��y�o�YҸ�3ƺ���N��x�x�u�]l�
H�'� m-�@�>�yޛ=�f�bM ]o�����O۲!���{�z���^v���{��[*Z�߼1_����X�rpIJ�x�?D�I��I���wܴ��ڿ@�pk�X�jٵ��_��1��*H�����������~�EDE���Fvz�*�yC��}4WQ����Ua���r�k�d��?qO�=�<�
��{�S:C�C ����_ղ�1���e}砋��e(ե���"�麿aC?Cǝuv�}���kY>g�Xm�`��hƘ�y�lk<��G3��`�+Y0�'���
/�	8ra��j��=�>��n�"��aK����5��T>m� ���D�6g�m��F��[���
��l�k 
�V:���3�^��(j�nr�?p{��fP���
G�R�����S��?�:�X��y�w�@�_�Y+"�^����2@��p� ��cA���$�Vm)����ET��6L�aJ�p�=�Oߩ�;�O�"��#������3��'�3������X���,�e8	N�����8��连J="��?�#�1+�p�q�������q�5κW>��2J�JO7�Ʃ2Q�&�D<<��
��^x�+PМl�zc��g�xI��)����t���T�;Q�9�& }O�sބs�Cj�T��o�.s��z�]r�
�����aH��ULE2�Ȑ�h	�e�!T��4L3����[Ŭ�6~�$���W���ǽq�y~F�7LA1g�%���n�MuNY[9����4���G��>zOy�G�Tİ���ǗT�Q���`$��� ���c�w�4�;�ۈ���N�(�D7��cr��-{,�4�-]�lX���q��4�7�d̴��d+d��1,ഃ�Ѕ=���7J��<}�S��,�'>_��䅲HP*w�5�1ݠ��$o�� ��i���3kG��DK�:��:e�q�o�����6��Q�3���놋�U�|���܀��b��ි1�aIQo�sm��79a��|�ቩ7"�K�NW3�*dĒ2���w�ld$���n�x;uzU$�+�[
&���@'�w;w��\���Ѽ��hWP!9FM���ul|)VHõ�����V��B�V*�e����h�;����_�P!H�α�j�5S2�4cӫj�����&�H@�l�a�x^y���cL� z���핝=��Pzȿ��u~�\�`-�#{@�[�:�ϲ��[ƀ���o�2iW���z'.�s�T��_��殚�=�/����u�1�NKڥ�Nx�_{D
�y9�2{��T�S9�-����b
iF�S~ݡ>s,��ݞ���C+�<?O|)�3�\�S�&��`���tc�ϝ����Lm�lrFu��(����yVN�M��ǑC�L ;D��r���+M���J�T�m�8=�Q��A ,��@@�����j��ڗ���	j� G���7&J��ľ!�rߟ�\���8A�L����-<"�_ݦB���	��{	�a��-�Z1�~�k���=cʥ#2�MO1�Z���w�2L��6D�d$�wI�R�%D�q�'B��P)��F~5��ҹo	Y$L� �'�L�B�	j�m�n)�l�Hӹwǂ6|��ܥ�J�?����S=���Z�F�on�W�<۞�#|�ᵖ����h��7ЂC�����=������H|C��8(|�l��&��\�#�{���c4{ᤰJȈDAdڠ*���|��w`��� �6R�ڦ�CJ�RA�7�Ps�;⠥u�=�)��mP��9��ѢmU��MQ�;��M �����c�%���K����\K���񴟙Z�������'�@~ ~@�!����E]�o�� &b��j�"k?b�M\p���5���9�z�}�E�.�#�Ō_j���y"����M�η�J��tY4�h	"(�^�R�טj
����d ,��/S��h �pFLlؓ,Aǟ��0��#5�OH����)���֪��{d�Rj*�+vӠY��&
�m�n�S��|����f����_x����⢢�i�Nb��LG�>Cm"�&l�5�������(�a&X�^H3��t���S!CԨg�E�����$S�Ʃ�v�L����I�ߑ��{��4�M�"i>zwz�W)��2.�S��$��3�H��(rX���^���*�*
GR+E�{��\4۬�cO1uO������I_!������U�ܧ)�7� 
����`�{�y��:t8��WS�i����_�sҮ
˴;@��p�[(�϶��)�Y�up0��Os�y��A ~�Fu|;\A �]��3E6��`�t�RN���ݗS���O(ᨗ���`�7Ю���)�
��ҹvu��$\�s|����g�ǃQ�X'�N�xQ)����$�����|#DGAx����3ϑ��b�J	��grf5}����!���bSa� ��v�8:��*�3㰦o�p��M�y�� \pr��pwa���S������k�(�(��`�nD��B`/iSS�f[�O���d�t:��7�9@��~�	����{��ZE������NŒY��ø�����_NL����\�|�Δ����s��Je��7���'��d��l>�M8��bܓO���M�55!"�I���dQX���]�-3����G�:����yz~e/&�ߞ9'a�/��Hh�
��N.�ўX%�0V�I8&hx�&D�ksXB< Imst8ctb�J\�l;=tX�c�����P�\əՖ.�#i+Hi}�E�@, �a��̜��
��Vg=��dMx��d�˺L.%���I�YIGlWcI�/��W���E��NC��xG҄<�����-��Y�`N=S.��&��}�z��y�x.L�Nܸ���3�>8��F�/?R�ղq_��
Uk�Q��a����fA
D�(M�9��z�e�v93�����(�n��% 4�Q�Y{%8��E���yD~{<���4݂~��kg���݅�m�O�c�q���Lc#�"��ѩh��>�����!0�9A}��m��f�c�b$�� �=�/���o�:ۆ���^aNҮ�g*f~h~�#��P���V'�G�Lm�ܸ��<m��Z�=��k4W���5v"Ζ���-!$��H�
�@/^+y�����`�id5|�� ݮ�6KG����%8�fn��7!*��[[cS����O�l��y&O5�R�DH�N�ڥ����4��(Z⌋Z�&tV�¾1�k��Uv�J�Z�����╫��������jt��4ZLoh�=��H鸜���ј��%$j!��
jѴ?�d��Y���+oဋ�7,�b�
5�
�Ԫ��k�Lн�U��M��!X&������a,�I��vȚ�ߠn��־6��K
��K�sj�}���G���D��F�p��.�W6�����	|97�W�#�6�	g����d�A��&�����1^�ˎ��5�>��'^�}J1��Ejb�[�{�l
k�����Uǒhf4�{�c�"E��Z�& �R`�ܾ,�+��
4q�:_�`��ۃ�ޢ�8�c ��5��+�''w݇�y;���!������,�K2w�����`B'�⿔Z��&�7������z��f㌧<.��Tg�Y�f��� �֭�̵E�}�&w/5������IbTK��h��+2��8S�/�Vo�s0�!�E�O`��E��"W"��s�UŕO-M�p��8�
y	_y��!�4���Y�GW��`%�.Q�$u�䚜�ӄ�l�77���`��3���J�k���a�۾������Tl䴄��ڐ%546$"�񸇝F��gn��ۓg�<E#�C:��b���*�-$t��W��{Ҫ�t�����)r�^u��z	l ﳌb�Qē�ucR��{�e%^W��x�9 �^�F�IL�����Z�ע������jn}Yƿ�)=�Y�M���VV����Bn�[i%n3n`+�ӈ%��t�	2�����q��\�A�;���(D�H[ji�c�Ɖ䠓<.y��|���{U˻�IÙ�r���KW@�X�p<��274�J,�VK�O(9�A����­ YT��9\*߼u��)v��!+�s��9��S�%�c�ƈ�|���]n�b��9q�C(5M�Ils9	�k��5��:��]!��
�C��=�Bu�sF�᫹�wR�Rf�:��0�:~���J'�Uz���)��\(}n,�2�QlZ:'��lo�y�`{��E�(���)%�G]�Kҏ��	���c��4��/�iW`w
a�?֯����}��GKVka<�'Ac����If�t_��$A�_*ߺy��l
��|�35*�U�����]�+��VJ� kE�����2�ƴ���e�O���K�w��w㑧ʲ41�劧�����`���<�����V�B��l�
q�(DAE�,+?#�����k��W^'&|�uA�@+�eB<�����lbN�)Q,T�!"�k��f;n�ߦ�d�xp��%~�c��E*��H�Y������ذ.���Y��f�@2?�*�uh㠢لu?���N���e��n��	_�UB(�O����=.�X��F}b��n��4���K��|���ꁊ���2����a�U�W|��z��G����\�[����p쫻#��n8`�&Y�`b��Pt>��'d:���{G%��$G�T�{x����+�6's�BG��(�3��R9'u�m=�C��B�����������ǚN���8��:ۚ�h�	������
���s2>b�J�F���W����,�zCS������(��e �bH����W�eH�����SF#��?���{�<�6�� ���wI�vɜgi%q���*@�M��A=HV��=9~_yWkQ�8�不aP���d0���3�<��%	��-^���B~Qn�f&�!l�m�.���o( %��p8�(jD�C��U�l�(&��Ko�nj��@���)|C����O��3a���P���Xd#��Y�Y[�jA�\���b?�fV�Qƛ)�Flk<g�!9Z����P�)�#.{�K���v�X��x%�%5�/���8E� ���#�c\T'��ygNh BWҵ�&{`f	��9|G�F j�;9{���<�)���#�E'�T?�;�����A��z�y�Nc]9��e ��粌�5�u�v�j ھQ��7�L�A����'��|�����o{D�6z��>���<sc9�?�	z+O���g��]|@�� >�.�I4s�\����q��T�3������@�kƒR��Q(ak��f;@c΍�5�N�d=Wƣ�l��ɴ�*�Q�?2�D_;)fV=��	<5-����2EU ��I�ޕc>�����Cz��BH�[�)$�O��Ί��}2n�.)UT�J��Ҳ����5����Y���[4OyZn9�t��H��(��TG��䙄/��Cg*!��W3-l�;�"���ۅ~�*���T#ʶ�dyk�x��TS~&�{��Q���m7 ��YU�+)��*�4Q���/��}PWH���>�y�mmط����}Sk��ݐVj1� ��+F)mș�S{����赾hC����m<6p�;?�ӑ`x�cO�%�*���{t%Y�N��zV@c���X�9Ľ�;��i�zЂ �> ڦ�zWʪ{�(�v5�wE�PN�t�Y4�'��^���D�ic��� a���@�s��VN����>K�d�:wZ	,�Y�1`>,�2A�i�k�h��XB���,R(-	O�/}Dp�6�x��ge���ق�;�����b���U&.K��\�	�^�z]��7Ԁ`jl���=K&[n�d4v����%Yyݯ�Ӛ�F�ޏ)`V�6��}9�Z��J�d��{�Δ��pp��������s�\٩m+k�h���g��p���6S�[\í���&*4���uu�����tB@�c�t��;�Br.c�$E�q��ii{V��2�D&�@#j��o8,\R���D�(w�Z�qkr��|��J4�hn
��2�~�� ��("7�9[�F�m�_�;l���@�s@R�(���J����ѳ�՜�H��<xM�}�\T_K��zqA"u(���ا`X�T�����X��\J�b�v��F\��������k@%ޑ����zٛB��qCH��x6Yt�i�^��9JL��~��;��6E�k����şxᛶ.ϨK�����ͭ`W.]s�GȲ�h��h��ښ.���m��<�|S�4a��Y��Ng������c�-�}svC!\`G#e(?Y�1Xoh&b���	o(	�Тt�p܄�PUd�L{�݆9̓�i��vX�H��:̧Ş�� ���Z�2��Ih8||��4	%�"�^�8e倡@�����6�`Z�2M��e��7iݛUd.������	6!m�~$f���� ��l��n�L�?<�O50`�E�&QVO����`(�
��-�����+����i���So��/�+d�a�	V����1]:����䡒F��R!��>m8!�<[⣑x/W�
�֢��5��Ea���2]��t��Хp��Jg��y�`�}���c��T�Z����V,��9b-±�L�x�9Jn�Sv�D�x�c�A8�*l?'�B�'���ն���W��d���{m���HwcZ� x���(��E;���!V���M��S�@�q��iv[�i$P�6��Z�+7Pn���~�Q}����c�h�K�~]w�kO��@����c����# (dn�@(�A:ln)F���+؍F���S�D���B(�������^�N�!S,��6����,��Z;}Ec��Sp���\������-��h[���I�� �j*�ՙ��lK�V��C���y9�V������=#+���8.E�캚ȇ�^p'2'|C\9�����yŖ�u'��Į'G�y�m[3�Kڴ�L|K �찧��B졀_m��2US7
ٖ��D�Y�_T�ՙq(D�@�pth�}`��.9��So��߬ECQ�UZ6�4	7�:z t�OU�4����q2����ݥ#������:�@�U���`7�O�j)O)�-$O�09�Y\=r���m�]l���k`ͯ�8>y��Z�@�s ����!���#���_O˫x��{0��S�s���Z�@@g���_�0�M���S��跽�Ljo����'�O�5+n�U�������FK�eI��L����uf�J\GbP�eSB�R��,�FF��C���h�6>�����<�+�6�"�R�sAr�ۀI���Q}���N}��+�1�4�^�3��pc���K�̒�l��������r�Q���N%&�^��,ϺE�(�8vW��hp�i�m�q�H1�g�5�Jc�HS5U ����{�uN�d.U[1��׽�q7�]N��F��BAD���/��0V����S�4�?%[�c�14��o�G�.xf�ML<l�}<����s�H2����;r�\�S��@jN�=�cg��h�p�TH� v3�sv�X�b{\��]�G�,�fr�eN=j���;X�jJpd!���t��c�5�t�<w�3��ԼۇF��ޭ�#�v���b[��=y5�`A�#��r��$�\w4-�z$�y�>@]��)]�jJR�XlxVHYEB    fa00    2e90� �|���X��],�M���C��Ы�_Z<9;`�~�,T�g���ȬC+F�Tb/R�K��*�B��Xi�Y�֢�ƻ�S�c���]{��HA�7j?���v�����A��-�Dx����;]���?l�B�49m�:\Q���WH`P�������I��n(H�x���O��J&+MH�jeX5%�@wD�:>vH�ȑ�,��ף���δ���:���_���D̛�轁)���9���g�����޴��Q�ekP���CCwG�B��BL�S�k�[��H�{
3p�Km��g������MnT�G��UG貘�Cs��� _����gF<��z��/��hH �F����6�!��?#'ykݦ����p�$g��K=%��>� �
Wrf��N�T=i�VA4m�w� u����9���E�B���(�h���z���l�y?�S�ET�H�g�ҧ�m��Ģ%���D�q�� {=���&�������l���9b`��(F	�������o���s� �0��+Q;���jwb����
��7����yL*m}�LԲ���8��"���+q�(u���(��bS����]�����ˏ��C���׫�,�U�,tc��p\�%�ྒ<i8���8�yŌI����Q�� 
�y��>�Ala�^�bA!�����]�H��`0�L@�ޕ2䫏�L�N�?$;4�����b�}8�v퓒p����`��_5b�|9N�Y�,aJ��Aj��ƶ�SNϣ1�z�����Y�Z4l݃F��w"�-�Za���a�R�o
��	��#[;�g ��ګV���"2����zF��#Y5��|^J\ǟ����v������D���-
*���v�Yfo�T�"u�,o���P���e�-[
�[(fu�J#�X�(hJ�x��i��D�����昗1OI�f߯΃�-%�rY4uϻW��P2���*�E�hdӜ�Q���5e�<|�b��	%x~�8���Q��8����-��#T/b'�@����u>l?��{x+�*p]����-SV�mR�z	��"��I��䲱uEdy{^i�2�	�� x��HK:�g�=����ζ�H̩�K!>�`�a��M�[��b�dH:G4[2����
q%O\���?h��G���O��k.6���+i��Cx�++M�۽Q��<��7�� ��(�i�˅�2[X;p�q[/<��B4������D��(u<���//��~�֦�82�Q.Ix?r�e�Q}�f?��QB[��)5ԩǕ�M?���;�n�ⱱ㣺KI���Vr�-`G�����ȋiث&E�~t1S���*�18 �4�pp����^h:=o-a&xZ=?�n#��8N�U���OF��h�v2I-��li���>B�J�b̻���-����AZz2)��w^�,v���%�w�c� ��i�En�ś|�h~���Hpٶ��P����``���g�����s����!�	_���'�:��_�<!(7z܋�Mr��d��$6����>�㭤l�]���_2Q��+:*���O��ߝ��]���	�bU(��������C^~t�g��`L+�>����T�T	!щ�,�5�E�����ġ�����d��������Z+Ua�Ua-{�:&K�/2�^!�J���3��������:�6��q^w0)�f8��6i�d��$f:ԫS���ߺzn�8nc��i&2�kXXV:3�;��@٘�s{��'��4�TL\(�V�g4�Lz!u&�jBc5�B��u�4:���_ɠ�dy��s�g�K-�y%�*�/�e���_��纜�ah��$�v\t�F��oSj�a�*U��ೕ��ҘI??�DK�Z���f���{��VJ�!��5/?Py�Ǡ���ԙ�W�����`a����
��0W[jP�L������ȥ���������� ��h���q�E��]Dm���(�A60�q\�l���1Yd�"��'� ��7b�����m10�.��2�n�$� �b�wC�֛	�h�'eg"��&�W����+{.1/5���]"���|�Ө[�baE��O�	6aG�]�%_"p�C5|�AP�	�`1M����N	����\~�Y���)J �ՙ������h-u<��Z���ĩ'��$ˮ�1���7��Q�=I�����-'�d�7[m�٥������0à�7�*1��Q6�%���;��;\O�y��$St4�S��܅��d�=^�h�9�h)�C��7+�Z��&� ���]L�*�4���N׈6����H�"����$���.3�.����GI��Y:���O�ŀ���E�\���*���P��m�u�a����N@͢���%x ��tȔbb��Au ��4p������ C��A��<7�J�@������o)�{������S��kޑ&�=��B�Ƴ4�^�a��]��?8�(+��'��%��H� �=�W>�	�N�tq���ќ����_(+�p������[|�����3�6��s�pad��	�ȶ�~���D�$�H`��&P�������GU��ׇ��^�o�/P���L���}C���%v���c:@�p�	$��8�8�k.����m��QZ���5e� �!���ɔ-m��I������I.||X��Z(�
ǴjS�B��oL����j)2�O��p��([�D�cM:��RyɂHq������2��-Y��d$b��O������K�M���YfC��z�+ۀ����ix�����яʩ��sF�d`��d2a'K(��n�b�@T�BL&h���\�`dB�t��( ��d�dI��)��ʸ��}b�CN�Ѐ9��/�^���}�gۦe�q٘7l�\GWQ2f�5�Ӯ ��7Cg�F��."9��r�Z�[�ݠ6æ'$&�ø8t<�����os~|��7����m����� Uw,(:J�ujb���S���o�Z�m���!j�����\��`�[L�j=ھ�&��n5!�^�O���<�Y�nvi�Y��l� Tk��5��o��F����V�uS�� (?��0� @6�~:���!n������s觊�`xR���ϐs�y,Q�������Qښ��T�\%y��.��<(b��ĔiH��]I�@Zk����$������!3K�I�8��g�;M�������7)L >� �<q�U�V��2��o,���Yt9AT6�V%�{<��"�
������ϰ;I����OkXH?,x����R���G�Qy���]��n8o�ff�&���+*����wE'L�S6��?j2I�W��бfo2<_)`w�uy�_�o�@�u�3�A�aFUzш��gٗ����0@w��;��$�WT��r�c�~  �+D���M��#�Ca*ɸo�,]�-��3����.��~ʎ�I�m{Q�@�9��i�&٤s�Jы��Dqo�`�E�9�0���M��E��46 e
�k��l�*!��Q�R��r�T%A����f��X�FX:̼�غ:sP)3���=��a���3���Zi����'; (z�~��
 �|h�Z�r��z�B�S �j���=S&�;�VT��]�Là�Ǚ8��56�<������UM���@ր� ͳ�����|KS��2����v��m5���Ͳщ��Bn����[��2R�4����-�
YV7Ue���A�T����DF^7w)Q����`"KK��re��5�I�@��K�'ꕵ���4-C-#NH|E0;����� $��?���;���u*�ljb��cۯR�s��ێ-x�2�X�L�.w3s+�RәL��+׌<�¨3j���O�|ξ�[]���j�[ł�Y�e�o&؄�V��k�~\`�~�׵���I7\���}1Gb�F��,�C͉%��CU诋�a� ���}�����f�6���(�N��*о�?*����pe���H�����W���&�ƙ�����M~L�w%�	7.!b	q>2�71�\����/���G�=����v���k���I`��B�c��7�NP�&�����V�Z6/�3ė�% %��[R�3bM<�ZZ�5��e��㳰2��+�M5�S��Z���I��T|� �g㶍;��!D�=9P��A����r�9QB�w���:���6I2�UUC�����L�[����P�As2���K�YWc���)Wz�Hq�A?HXǀ�`���F�a-N���U��\1�����LW-|�rY΁%�T��a�`m��H@$Y���%®x���G�z�N'�i������5@��l�A���D�ܭ���BƔI���R��i�b�g.�@]:��ZY��@��l�	!��hǁ�/"�}�k�B��8ՠB��RMN�)�39qˇֿ�*f�g���p��7L�Ɵ�]�v�P�v��5��u�����T ��)=3�Ą���k	����:ȂE>�]a-��H�%[�fh/
�Gk:�Gi���GB?2@T;�����^>�����'������X��Ȥ�}�&�A�˲�Q�{������\�X��J���Zo�I�0#�ebp���B�2�Ĩ7���b�����fJEeIvF;2ґ�VE�p|��b/^�1��L
�UP5v���We>��w����F��/�])J��"u�+j�B�G�&����O�Ͱ��f/1=#��x�F�4q���d����!��zVDCR$�d݌�"t��Ov)��*�3+���e����)�%T��fm�LV8�cAG>�y��
J�%r��g�?@�Z�0��F�.)&$� 6�-��ũc�MɴRh��7��#`H�t�sY܅�t-hFT!_�1��9�T"���/��3���G�?il�1�Y����Ϙ����ǻf�P���%�����c��I4LEGl�.�}8O� E���BX���O}ҵ��EcI�+) �(��5�~��·L}I����ds��y�i�\���r�_�;[B���o��H��҇"uH�K�.��L��s k��B9-h��_�V��IԖ��z�yԅk���;��95�ƹ��I�#�^��3K+Uu���|f��>p�!�����#hgDn�g7{Vr�`.䨓TJ�1�~aezVy:���ҭqB�kqM1'�����<x��/�4ڠQI���<�({��!i?��P.��-Xz�	�^��j't�Am԰����j�qau�uoS�v"�D�%�eڈ��,�[Q��5�.7�^��x:��֝��Ȳ]"�]�HFjs��s�S��n�yQَ'�-ɐ��O)��1���+`m�틞5Z�����g�D3SE�w9�PF�]�ua^�x(�gc��6�8�G�˚���3Iu3J��̻�s��X?�&=��x�$�p*��w1��e��ZLOm[����=���Z(H�۔8��N5uO{��J��LW�.�� >�R=�A�ʙ=���0��.�_�<��U�z(�:�:7��DcEo�h�(OCc�G7�`U$��y�������m�p�\P��2-�
$��LX�|�KPys�(o���e?���/}|��20�OD��Uf�vY4A[��a�I��'@O�p"ʴ��r�>��ƭ�Al�@��w?J����Pu�<��@�7���g��ɢN�j�"���)���p�t*��ˤ	��>S���!�!M���|�#>Tq�3To6�ev�Y˚A����4���$[Θ2S��Q�h���ہ� ���=ao�d<M:��(�h�қpj��L���@'@�n�/��+a�� ڶu´_�������P��5�������A�*=��O�v��K[��8�X�'�݃�n�Ž��̠�lC�
0 J���Uz��͜�Y����L��ӏ	�V�W�r�E��K� <B_��6�v��u�=N}���C*Wc-�ԃq4�ID�ym�i�7���{�]���ң��"�B������\���\�jgX0�Շ~M@ĳr� A%dSs�j�j��1�4�Y���GZ���8*p��4�ehΜ�*wqf��r�*Jmt�����#� _#�J9`bH6]q�a��$���
�Sa�ɢm��:b�f��z(�??P=y$'�be���r�ox�Z$����1�㻘KlG�PK�/<�_�BT'��`|�����tN�J�^J,Q*����B]�o��2#\zLi �"#N`#���t��yb�y��Hr�@��*�?m۳��D��k.���Mȥ�p��k/:e��"�"�}`#���(?�o�o�@a
1���_8�3Ȼ�<S㌯�6�i�E95�(w"�0�����!�@;>[��q�	O�i�`����Ս�l����$�,\�Ϡ�1a�aq��/�)t1����
�c�����B�ٻ�_^�aͥ+C ��t_Tg�sX�Q�Ž���U��݉
�K?�apֲK�؜sa��S�9Z�*KvVy,x䮏��M��+:�G�9��{���]�?pl�#��R�̭�J+����O���wc��j�isΑ�I���
e�/o|z?���:V�ޠ��WB�~�����Z�R�dT�0l�z���~Y��BY}M]V��e���ːf�}�o^2�D�	�	����� k�4niyr�DcG�r���fgɑ���`/�?�ߒ�Ww�����륱�@�>�ڡz�E�ͽ�b
�;���n�����:���֒�7�S5��E����(�v�JgV<o����dv�� 	�'�P;5A���� ���b�ֳ߳��W�2x�J�s���֎��Hv`*+�ISi<N�= �p��K!��OǞe�,��2��6�$+��*��k�U��QO�W�O3W%���T�ը��0�׎.Oȯ���`$Մ��̩��3v�J�:����8��v"0��F�Yj�έ�S�� #��F���D��ڦM�2PV�T~��S׊ q'�*�
�*�&�-pHG��>�>�΀�b.�0�Y���n�xGc��^S��U)��H7��PVT��/��S�{�iU��W��~3i��Eja-2�L�0��*3���Ƅ���a�-ۗ�_��O�m�ڵ�V¼�7/�`�&���=��V���A%le�
v��ۭr_�8��tϹ� W�o�TL
���R�$E7%&{[�S��/�:�PAt�ʁ�D����f���k���p�.�`���EP��Tj�{���LC�j��9t�f�9����=��H�}Q���>�1��u$�6650��4t=�]��*�1��;C��G�D4E�g_w�h��u[B�{v��h�g
�e��rl�g7����<NL,(D%�VE��)�$Qo_u��r<����9��uH
,�H�2%F������(k�u�{9�=�?t��#Q��g�,Q�f�'�˦��>�.F=�^�-���<RJ��xp�X��׋x����ֹ�������r0���DL��h@�V�)���!J�}Xr�j�l�09�5���5-�z�{5��=��6����U�_*nC���_���~�\S��Dd���K%�+�>�q�<�;��7�U�O��N�����Ӫ��%��[��=4K�I�����"zd���w�-��L�m��p3?f>:�Ò����9&�/�����B#�^h&0̵$F8U��&hfdw�$rmՍ�>}�xzʻzS��"Mʓ ���Cwm�6o	�H��J���|�xE���#Hަ��ڴJ9,��9������m�ZI����<vR��M7s��:�B��4�=�{d+DǏ�2E�=,�%�3������w�Hv�V�@�`�U#����lFz���ʰtos\�׫�^�Wd/x�r헀��zi��|�$5���~�Q��F#uL�2ﹴodF�o�B�"̗��2�wQ"�?�`�oxT�6c3��]#�H��pDyN?��v��д��!-�C���h�*רF�O�#q�������7��$���ņ�BI+�!S @�G���^��U�I$��xY�Ll�y��#W��Ŕ#V�g�vID��@|�T'���h��C�x|N�=d�!-�Y����͊��A,ϯ���������qf����؆�!�"=���起��
����$��P��^g7�X&��Y�S:�˰Im��!H�V���~�8;C�4 ԕ���o�E�A�豻��T��=�.����Q_��I�e�NE�~3�X�)�`����A=��s u��$QUK�7O"�;�X�i�0���;�n����%�FXf^0��|�g���"��5!a!3W�����i�Ԧ��sv�B?�l-|g-[�-��1����l~���	B.�	��c� L�7��50��"�*{��M鰮�mD�*�b��.[v�XU�~����_��1�4�㶄B"����x�j�'���0���2�F([CM-+,/�c���X��GA�9?�� 0ݵ�=r.&�{�uyu���Y4�B�%�75r��Ѹ�:*��i̪�Z�qanã�����#Vq�&�IJ�K�Hԩ<�]�g�[�騣�9xV��OL�DQ��u�#�$�$l�}��%~��!��0��૕i��V\��k/�6&��NOەgHt�hT8�|����1*���־�x�u"�c���_��*D��5�NS��+��C'��=��s$]���t-xH���8�94�A�&��!�yz^�6W]Ѥ΋O%�ƞ!0��'!��e�\�<N�d�gD�n�[�����J��#�wi���Q�������d�����7�t���9��VX�WWXAc輻~�~��R����`�[���i��7̍�r�R�^�洔��E<��	:-�d9q�BG�e1��έ]B]����M����<��:}'����;�M��B.4DCT�������5v��J���Ӕ������&�����'+e��ծ�~�����	a�,<]�ۜ@�o���tSئ��o��	���`̷q�1jU�}����נ�*�KsUC]>�� �xKq+S�����吿�I�Ց�w&��2�*+�h?��F�;ϵ���q9�;s��o9���j=����w���HL-�([�Nߏ�þ��g�g��	+�Ӗ9A�ߨ'�e�
�O騟~�Q�I���9\S���E�"��� I~Q�Ȫ���#u���|Y���}��DJv�V��j��S�$��MA
2k3�Xad�
^�4���hs�Nʳ\��ox��l$,��]l
�;i�=l�{4у
��'ӊȌ(=�kؓg�ҁ��y��a�V��s�s�e��L�.@	E	m�I�����x��2:�|��_�q�ey�f������ɤ��(|1��GO� p�T[�&)�n#��S���6vS� `jT�k3U>���¡3�k�@8���k?��ĺ���2O������F���>v]��4��>1���'7�Q����)Y���t�U�$�������z}3�w�_��Hk���f`@�7e뷩U���P�;�n�a�n?1��^E���T��'�.��T,	�p0�:�ҽ�?*M��/g�J���{�%�Z�Mi�����~����"Ϸ��Ѓ��r�Q3a`�JSo�I��#|g%��b��kpRc*����K=����4���Pި��K��]$�?�,��e<]"Ń�ǆ�|�:$#H�wG~s!P�¿O��HBI��E�iĜ�A-�I�Lma����i�X�2�16�DWC�r
y�:���S���h-����L$A��M�����zC{ˋ�Z�	�\���V(¸�V��)���������&�2�$g��6�f�yQ���'�!�R���f��Qω(.H�6��ia�G��T@~��ck��
��e���.��� 9���o�o���*���f?����1t���Ӌ���]\���x�~d�����*�8�MU� k]Jčg%g�lWi�]�o2T��ǆ��6G��b�\X;�ߣ�w�n��+��<dM�a{��'[ڇ��T.N �����`o���)����{�d��-�H���U��z�A<rU���V��3�^�n����0���d*��_o;l
6�G�q�U�q��XrE��*��g6]j�	Ѽz2ʴ#������I[B�Ŗ���|F&��.U����}e�=9]�#�N5W�#�Ь�ɍl�Q7F�V������c��� �W5p�qQ�y���­!�#Z��SJ������8ecr��º�ņ< ��`�AgE�a���q�P���Jb�,(2s����o��aK�ͪ8 �aǩ�'�&���F��?K���"��c�r:]սY�u��yF��0�`����(��&�2D�W�*h��7�u�/�wX��r*��٣�u���LvkG�D�H�ـ"}ks�%x����zT���9����gdU���A����uB%�(3���6MY�����yBXx+�e��S�x�&�@�m��s�c�g�a��c����cw�)�D��}�1D~+Ӆ�$E��s�f�����5Xb0���e)V�i0�TQ���5L�̔d;D��%���G��q�ƾ36�pA��l�Rn�V����}��d��-Pƽ�t�D����ص��&f*�%a�=�PM���c-7O�ew�o}���Ko�+e}���?�y�4l���T���*�G�t������Nk����?X��78oB�Ё��������`M�j�Y% 5}$y�_kr��]aV�����h�f��h#�����К�)��"���S+�Zp�*�S�r�Wdv���H�?�e�ƺ�Σ�N���yH^*��@�4�
Y�G�ħ�$�+�6�`� �aݚh�t>��C�iu��6�ݪ�zA�zwe��d�[$&($�<;����I���0�8���Z�A�+'��>��AZ��ƍ!��OP��!u��v������'�`���s�*�S�|�/�cT��W��zQ�:n��l�Ud���)F�P�����7��s��e�ֱ"��R�:v�(�]D�QÆlG�j*��?�5�"l�)za(�;@�ݽ(�3.��~TUV�"N�&�����3-@K>�������GBk����ut��[��u��M;$�It5p�PH���v9��+9DEA�S׵	�)� ����t�Q�+�T��N[�K��󘗗`��QC���񰕲�yC"�͉dчb��CMx��k��������
;?q��¿�4��<b��79��]�0���c&t CԚ�}�!���B���8!��âFQ0*�;E�����s���_���^��ܯ�-��i�����h3~��
c���s#t|�jQ_��� ��ԟ�� ���r#����lQ�[?���[�D=m��V�e��.��3'�E�]�fT�&�ݓm�К�����|R��S�p����R�&(W��d�͎�C6N;�`��j4�b �M��A�}�L"ʹ.~Zl���dn�!�Z���f�9�'kЛu��Z9�a�K5�M�Z}�:9
�קzL�i�S�+�jt'��}��g��`���B�o�g㩤��۶x�I��K#����Mj��@V5
衔�-֔^Y�����Nc[�aԧ
��@I?�;��T���B�$W$�6����,@�-����{�uDǶ��l6��np��'�79*����hZ��j{�X���":X�\SqJ�2��p`���&�r�"����7踊�l�ᄺW������Q�e{Ddȝ�Œ~��y�,��2�7;��>0����mAW)��7P��T쎁�Uؙm�����:�o8�
� ;g18ћ�����7BK��y�z���|��|��!U&{U��a*�2>#CQD��G'� /�9oyO���K�A����\,��Nz�� ���=���dK
�-���!XlxVHYEB    9e01    1c00�s�w�jv�c��B�:�^�lfF����V:�Fg}Z�
��f�7�'c��ڋL�����Wm$�$,��fq�W���-�j�����X���8��Pf�t�L��]ba�5��x����Ŵ��?��T�*u�%"q�L�inn�	`ed˙��K���|`NŢI(>��;��(�nϖ�����^����+&�o������%�d��Y�h�q4�����^jz����Mm�C_8��'�G��;�p�; �K��^�l��7���n8-�DZ��x�AIn���xX
cf;�����)U��3E�ق1ݟR��hI�dX�[��'9�_!�O7�a� r�o���J��5��7PVW�ΜRQs$\4��3������P"�4�Rj�f.�`��#��^�遶F�pV��q�`��I�9��v^	__ս�>�rA;L=��Dk�j���k��F�A�<�MQ豋5Y�r��5d{t���٤* �Ҭ��U���r7��{��}�O������b�S���ʯ
�2g�����x#r�����5`,�q��X@���:ߘL���5M|yiE�("��q��3_`�0AO���Vv��$��-�����A#���d� �P������q��t*^���,��-�nf��D�<3A��+%�䐖(�;^�;�1��Cw����>����i��\�v�%c�k�6s�> �]����bSR�hh0���&��v�e@���fl��=@l�irZ�'v�z��Q�2-��p|Cz��O��;�M%7�uh�;tU�t�r6X��ğk,S����A;��B�8.P(�=���k8�`�&����@x.��a$=:M�Um
@P`H �y�f�5�NH��}U1���Ŋ��uj�ocp�57*q�tw�%�)e5X:欩S�i�'/�v�<�=��=��Y�ju���D�
�P�7��f}��x��>tī����h���"�q���@
������a�8i1κ�@Cv5�
��&(f��^�Y��N%e��<GNX��  w��0�F��4S��j�ГUa�=�'��#E�w�Z�X�V��U��:�W|z�6}�͞��t��A�WH��S�`NG"[��K�N�U�����[O����W�]��W������R��V�@�&�<s�K;dITƩ[�|���-u���j�ʇl��t � �50�=d���SL���쿪�QC�m�^�~_�/��/��R�-c`�$�������	���ֆ��U����b�i���r�)��S]L�ԓ��@>]K���@���A1�;�LE�(�+	,�=ĵ����H�f!*߮�\mjx�
�VV��/6)���$�<���s-̀a��C쾗���G�2��.���^#�0��,�:���ue�KM�\ �����4&�'	i��j�.��e<>��&- �m5�N���lPC%�_)'J]P�6�)���ގ��w��ˉ���8&{�(���+�Aad!	#0�P����/��%����p�6[=J��H�����,�vP"V`���@�ecJͩsG~�BĶ�W�'����ga�2�:��9f�:%w�WB�H�C1��p�M�f�i�[��D�ֲx�J54�SFr�ٗ��F� F�юm��c=��=��]�r�H��])a�b��ReP�&8bh��,����,���A[׌Y��y���`�]<N5חQ���'�,o���L�5s����9�Pl��8_�Q�Q*-����xɊ:BA{���v$�\�RC��Cl,�h�c��9�j�S�������ɷ"�l�����|n C�idՉ%��eM�� �&L�������ޫn������m�������i���=�J��zD�kܷ-f���޽�2+^��-��\a���L�FY�[���Q,�*fz�C�T0<��eZ�r��3Co��?��7����9��~P��rD��XY�/���c�8�X�?B�m�~-@���*^Ab�����|�U�)��:������n�`݁|�S�A�E �5-��^	y���1Y���N�ݰi����_&W���1J`I9�6#�����&�lRJ��%�(F�i`h�_�����u#�3L>�A�cL��A� �86L^��(:?5�9���n�mR�B��f�q�teo-6_8\��΋n��LĿR���#�R����Y�UJ�x<,�aBk��B�W�X�S� G*�� �TMrr!�N��0�j:]y��]]�9��3-�:J��<s8��{���Ǩ�(�V�,����tߏ��,K�cEW��9%p[c�l�I���&�,x<q�J?��P�E���%�2p��tR"��Ш�S�̫6��ڐ̆�W��'���+���w-� �兂ѣ����8����0�0^Y|�on���%��lE�ɘ�рgڌ�ӵG
�.߉\,&�Z�3j�ֽҠ+S7ߛ����|#�EKTD6 (�p�D���n箬+�&X��#N��`z�怠qԢ�e���q������hщ�wf0�^?��}�Hr�Ð^��Y�������>��׵��yjj��fv�,w9�� Vt�[��l�ۡ,��[�E�����W�Q��2 <�{�]����%��D7CO�~��4�FMn-Ϧ���ߞ_�Kv�x�2:����R��8V���4 ؀�8?@�HHT���b_��:5-��j����A���@S �n����X����ۡ���~���\���6&�(m,3��	.ā#^�t��9<�[�Jq�t�_]?∗H�W��D}\;�����&�߼�Q@���\���\��^G��j���5�����g�<��k�Z�M��=K�����fV��X�Sr���n~N_�㔩>�����
�����K�|3/�[0;.��m�6�]G�B�>H��[&��fMX���cu�[���LU��̛-H��M���pyZ+$�K�N~lg'�?��r�';n.JՓ����Ă�<���?��ٿn����5�L]��O�����^8��4^w�n6�K��6fUn�N���-�'���n�*UI��+{Ž� ��CE��o��38�{>uexq��cMӮ�-�!�y^
 �k��T�c5�W��T��>�rW3��O}��35�a�X�<��f��h�����6���6��e΀�H���S�C�DX*c5�=�}�g�a�M�YPy_��F&i��Ƣ/Ʀ�u�*�BܜGR��s�����],�~ñ�a� �"r�D��ؔu�����rr/����>P*l_U�1��q{d�o+t]�\q�r��)w	��߬��^e6G�AL���CT��$j�1H�[h���7��-\�!@qg)�UH9�ǅ+���f$�QM���nډ"��+"��e��@\W�mtS�  ������>/W"^EQ� �v^�&\{5�t�q�t�k��O�����j»V�(��w�mT��8xW,��HT!����l�VY�	��҉DtĶ�m�]	���?w�,�Uq_Koo��(��$�x\�kn�O ����ʼ���*���Y�Ғ.J�B�(9�K���˷�ʭ�a��0�����/Mo a���P�+*����"�m�����	��;����P7mZY�a�Z&Ί��3}�7,��]���"�W�깢�Ǹn8�M�E�'�?�H���2�
���QFV�t�.x�7d\�[������٩�t�׈i0�C�eۋ�~�y@�<�����NpRі�/��T���1s�N�A�פ�ɭ/��5�vS�T9ʰ�m_�n.noN��-�k��w��'�Q��B���zr~��՗
����O�&�Gч�!���/�:ػ�Su[�u�k�	��\p�U��mb-�]ߞ��ҹ/(����B�^��b�`8��8-�/] ����z�m���6���FLx? �҄���38�{+J�(E�	t���4yx���=Z�P+`��͔���K.��g��j K�}ڧ,�q��`jl��)����c�ۗ���
���q�5\���4�Z��1����fx��]rG�av��$�J�}bN'�����\�[]b�P�c�]���-��������Oca�B|���!�Y�r����9����aC��z�~���"����p�9A$��W��Y+�\�=;���k	�d����z���aD�����[����M�;���s��l.�ܢ����V�-YP��'NF����YZ������ㅢ����t�BEi�a�I���q �aO���W>h5�4!\{�?jK-Wi9�j�g�^_�F�����^0��r�oYN�b!"m9Es�o	�]0h�֣.ͭ�!)��ҳ�p�bZ�n+�*�	}��D�Vxּ����d'�=�*�����	(����0�K���#�������*��$�8�����Cst#	�WdU�O��
(��Q�����jQfՐY#���4m+ݕ�M��d
�5���¸1�d��⨔�į�]i~kȶM�K����١o_�S�Sܬpv����R��{���(��Q�f�7/���Z��o��h�"��Ue�*��0N�}O��><�y c�i�5�녴� �DDː�}�E0��$�8���P+�S�nR�f�Z� �Ҡ����s_8[x5�I�I���"c�b�=}�*�>�$'Gl���eũN%�,��I�' �]�to�Q��咧7��4ٷ1�jx:����ǚg*Ч"��#�f.������Sro��or�m�A�ދ
z��7�{��y&Ԉt��e�0����%���7��܀Z�|�h%-2�T��o��8�t�.�@K�oa�����\^<�O��eA��򷧂�p��#c��I���F5걀��jX���g����~��.I��IU<z�P欬�)�F��+r��л�m��n��H��"锘�t�d|�MHʛ�u�p5��(^�+ );�����lV���8��T WP	bCc�$+����.L(S�얕�W�vjD�?�E+�e4������@�0h��!l�ԩ_\�H�@��7�*���O��c���a�&��d��V� ��Ե,z�W��g�oem9:~�w�H�-ˍ�⥚�1�ǩ1V�ΰ�Pq֟8¸f�&x	�(����_��%����N���<-�����l�$W5%�er������W�t���j��z4,�S�t�"S�t�n*��U��q��f�>�\R��;����⁆����5��$�J���`�)�G��=:�2D8;��]�|�M����j�9�]��:Ҥ�^��{)ϫ!��@>̼m�&���ږ�e����f _����M9���P����^��A83`Ƚ:AVGT �ꋻti��v/���]*��Ɉ��U�w8c$�cY��D���!�#�5�]����3����?+��[Mj��=><��)��=:�Oi�ޤ�����~Q�4sW����b�YM���������7u\|���]|�?Bbe��5B3�=��\P�|{&�Ej��6�y�T9�� !C�x��R_�I��?��j/B��҂D1U�w����n"�|�H1�k?۴`��{�����}�KR���Բqz=4��,�X��Pw=�_Sf��fG�/>v���������t{��*+�ц�l�EY��&�P�W\���fGޘ��#t�l"ޗ�ʒ���N�j���r�=� LҸ�hMu�4�FM���/<����̫���Co28�7G��e�=�T��͍ ���ܲr�C���Xֹ�Ub�� K�I�����ڇr,��}[E)����Κj~���J^!u;�A��� ��8�<�^��B�L�/x�*H6���`����O��DGgt�X�zH����hPm5�t��+��nS��K9����d |�51�0+�T~���/����$��l�������+O�2?Cw�~d�ĕ� � ������lM��D���Վ�B�@�8�}��&��vM��4?�E��Չ����Q���|�ݵk�8�}���ˏ����n�79^��o��:d���j�J��.@��2e;�� �!Q�2/³�f����s
d�h�E�2�eya� ���/0�<�4'���%��
z�C5�69�bظ
�(�;�f[T����������l �%�qRW˕Vќܪl��&Po^��B	,�k�PӺ,��e��m��Ɑ�W��4����(C1�$��#�+8@�������yv����㯝H3ۻ���
]6��h���C��e��),o?v' ����B�2��������{��r�F$V�\��v	v"��1�Dk�����B��29�î���~���ϑrS,o��?��3�6A�M�����f���[fP�u�o�B�����âv�^ӅЙ�#�Ć�cՎ���,���T����t�$?6�~u���'	���c��m�P~Q=��H	�Ճ�����m���S�ɹG����=�YPHt]=�����eVH�LN�(�o��O��e㢏�I.J�O{k�g�Nj<ѯ|E�2�!&G�]_�/�2�����:'�;�su6�?�Bt�u��V�K��S9P;ɋ�}k��Һ��'���iݼ�hI�i�a\���Yfџ�&Q.R �g�m����=��Ůh2� ƻL��S��B*څ�Z�ݲ���\�~fm�tc�ȝ�.�{d�b��t���B����O.��q$�u�R��[`O���	�
���
����1&�؁�Ӭ����%U&d�H.��~0��(��� 	>\����3&�;B�V��H�)�a
 �����x�n�^�&ͧS��!���ha8(�%�hx% jO��2ti���o���!]�/�A� b�0����
6M�NV�igx�_��_1. �9���H�I����jGc���{�1��(�v0Skn�}Ab�L�̂Ћ4�h�����&%�X����N�'��Ɍĩ�톧�����>g�Fx�,.������ڴ_RT`����j���x��8Z{��d@��+�%��#ִ����|���[�m1X�5s�������ҽ�FKE�k�i��.�1�A>���ܟm��2��I�i�� -N]�d�����+i�1��T�}�?`*f�_��tR�/��;k�n�_���p݀��-+