XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���^=�����s���Y;������^gOw���[=��k�[{RϠW��mOg�}��
<z��渿�+�b-&Bh�d���K5"���	��S�,%� h	�i`�i�kR��w�t�a�����������3�� )��Q�t٩�D���H��
��!s�r�_�V]�n!�|������~
��]��\Z�6Xr}��#���쳡���υD7�;]'ƭ�1Cb�X�}��6k�^ڶYS���۬.2tl?�X}�
����`Q��(��U��
-��O�Q�.e�Y���ӫDS�n��`�F{�w0q0o1\��'�#��K��3e,jDO��P�\�;�\7�@#7��'uj L�}�4WB,�}̓��g��c�燾O�Ru�`���l�{��Brt�B��RK��n{y�1�bh��?/�<F�K+�T��~����Rͺk��P���,�'@wx}�q"��%����Ѹs5�,��+��{�W�,�3pVF�ne���?��]~��ɗ��T�C"O3 �1��%��}�6�\��sJ_�u�~���IȦ[����q}�H��DuF�u'���.
����_p��tj���ˢP�¼I�;WűU��y���P-Y+���|C"e��|����N:�6	D�i9_����Q��<&�Or����S]��g`�j������0J�����l�Ue�+B��[�ͅ�O拧�m}�#Z���f�I�����":�<�v�:���+��]�WXlxVHYEB    3ab7    1040+h-�QF�q�9�f=��
��r�y��FM���hC5%�ņ��<�����a�j*�4�*��M6E�?:u��^�	���7�Жv᪘WE�n�������D>�!ۮ���I���Ws�e0�6�^ e}���fӳ�53�
���ͥ~.p����:#��'YPv���m+z�fDQdpY]��*|��g�/PIJ�b�Z���7E3C�u1��W!�:�,��E�o�Ef�հg{@Z�XR.m�F��'z_�]���}���������Z1��S���oC�4�li!<�S��=D�b<HT{�΍,z}���emS@�Wg��a���c�f����0�d�j�ͲV�����E �R_����b˧~1����8��x�w�΢�x^~��N�G`�Nj�oU�k�q9��o3���A��k}�"�LD�|�E����������QF_t�����"+O�gm��ډ��t��ҳ�n/�<ªW
�,����8����d�/�3K�y�?��U�/: �m�ҵ*a��O}�N�n������IAGs�2����]�8g˙�	��ҷ�I5�^��������,�jXc��D?��6s�BS�t�+��@�*��E.��I�'I���=GnϹы�Q�7� z����b�
G����v�52V�%e7>��&��;Ϡ���[i#����r�%	c_�v���@��+���ꊢ�H�Ws�.D��)��������?ii�\�_�����@*�������U2vx�&"@&���m<��^�V�r�#b���nt���߻4�*{�#Okz?�U�Ib��S*��.4��
��k&.�mf1�zOd22�MGj�[��)+��}TBt�mZ�"?���S���l�nU�*x�P�I�s ����A���r�����u�M�X�3�8��,�����
�+&��ސ2�[��Y���7٫w�q�^�(��9e@G�^���n�AF���PjBd^��cW-�m�ĕXul��"a�P�z*;�o&%��9�t����
6�I1�"g���^ֹi�A�i۔�gd����Ê?�AMZR����X�"�,/zo}��\wLM�W�e�Z6ou0�g��z�L��%z"�{֗˱6y�m���/� �<@=
�u�L��hh��N�J�(Z����j)���ɧ� ��^b�OXW(�.[i �{�KqA���ŵ尌A԰���:�/F�Ҝ����Je����2.4ݩX���v/��Z���Q`�i��&��e���58�2�}��)��j?���;�D,(:;,�Q��S&�^�5�2M��W�,x]�l�����4h�'��H�U~��"˒�,ց��v���\|�fp�lg���.����TO�u J���k��2=�����؞ꦕ�w��	�M�>���V �x}l�t۹N�.�J��A�Qo+�	6�Y����@�8e�Ą�8�2�t�@ŏ/,J�т�c���k��_݌A	���ъ��E�~� ���5��8��k��)|d�V6��/)0.̌120C����y�rx���$w�b)6�k�ZvZ�ʎ2�}�Cyy�ާ:�C{��
����~d���C�Wi��M�&�N=�n�w�Qx�4a�Q
�C��:>��^ Z-����k!�[�O�]���D�	��FH�
C~�ͽݏ3���6	�%�<��!x�X��o�,�`ʟ*�r�#��?���b]iVg��.��n�L��V������6O��B�k�}l^��|������Ss�� _[�9g>��CBv��ZU�(��	ě�!��G���/�jk'�n=v�A6��`�;*� e��\�`/�|_�u%!nʈ��n�D���綒�g5�$!!�	}�ٽ�wS/�Ѫ&U��}��'�b��E������ύ���;��,��ۏa*ȷPc���DkmA#�]"�m���Q��8x�y�w�ˉ4���
���N�	cTQ�����H~���� b)�Ȅ)b�6�A2]Xi�*
>�DS�?���9v9T�F�O�k�T�̲�x`���6	�b���g���!%3OS�&Z�բX��h��85`	%��AbXV؈��g��국��c*a��sH��-Ek�Li<�Z��uӏE5n߾A�w� $���}���,J�-Ӌ>�Jšrz�u,o�)�v�E��Z�ݧ�=@�</7܎>zI�T��/�dJK�`��2��c��\��Z�aQ�m<�g.��� �s?�����N�qsx�"b�����U����ې,:�*;�Y+c�)Ly2gL��Ɍ�KH�$],��S~�6o����գe��m��cԘ�q;)���-�Y�0�V�gZ:�C���F�R�t��&���W) �|c���Y-.���H[m~�oT9. �\n��	L1�EA&�p��}�0s�&=��i7�G���M\2��/~�4�1���%I��S�\rEG�6��t�u!A��[Ɏu�yHw,�i��9�ˁ����_�B����DH��ۈ}!W�����!��ș� j�?Y-�m��>���Y(I%��=� ���T�I�!B\���e�`�Lw�K�9�gY5��P	1Ua��Z���sI��"�"�X�p|-2$t7�P��!�MMk.&�3�V���:�_�D�M�hﴷi����-^�u�(IX�LP�V^4~O�i�Aw�"�U�Hݰ�Ɔ!����j@b�����0�!~��(�8���[�2g �n8S�=4ͻT�p��P3q�F�O]�S��k��X�t��ͳ�wO�nE�D�iH��p�JIS���	�V<��;Hz�Ӗ���g��g�n-��G1������ �r����Fw^!�i��8�~ş;Z���@����\'����z��.��1 P�4�ht�KQǒ��Z� 9����./<����N�A<�{�ֈ��Yʅ�.����X�.NбY>d��m��x��4e=	��-f�NA*:gR��[��0�W�+�wm��q��['uq}Fd�8�����y�����
_�o�k����mbn�dh���E���ߵ`�(V�r�@>�Y��i8�X�ew��WM'��Te���6U��Zt�e��%���4'�]��(�0V<:���r�{���w�G03��47{�B�n�C�vuO���{3�w��S/�7h��|?���wm�N�wل���Uub�8�
m�|�=r���qZ
 ���Y`hl�	�g�RL�׉ jSɬ倡Zӧ�(Gզ}���;����o�z���o��׾�� ���q���!���2P������KU'��m
�BX9c�Fl���ܫc�"��Q�,V��aS޶\�&�h�
4� Py4� ����[�����-B�Cu�7�F�~���p \ �+o�k�v4����y��RS���rr%�X�rފ�c�U2���s�#&DP���L�'���)J�G�Y�o�ԡN�V�IWw?�Dl�LAЋ�1N�⚖�,��'�{DL̟e����K/n��.���b�Mޗ۾
م�l��:οDm�����;?�R�TΔ�<+��gB�eo��O�(�%���^��0y����-��+�B/��S���N3�	);l��a)���r�	?���"�t=h��m���Y�ǡ^>6�\Q"�*���FN��'r�,��%"���ղv	Jb��5ډ<���밳�JO���uߟ���ŅQT��K���he_3h�X��ŊQ�ȝ��{H���r� �셄��{s�Y���SN�t�C�+;o���� ?���3�ĻEv3Pcp���nn�F�S[��ב���q�OF}��b�n4I�`J�m�á��M �k���Gf���	�9�q?q����{U=�UAͺ���M=����Ź!��ߟ�{l!}W�5Ӕ��P�؀VUo�X��'�X(���,;��|�_`�6���@��."8M�E�9*�:����(�b�E�Ǐ�����11JW����{~���MހU�aav���1�=���Ӊ%�w_'�B=��~(��w#jS��\�%��_����%zP����d��0YWp�}����)����.�MT;v�� {�`-�-��I�sc�s�>��v+��1APz�����)Uahr