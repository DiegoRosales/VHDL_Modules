XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��d��I�g^겵z�,X����@H�#\,�mx�����gh6���#��A��u�ޤ�r�ߤ3Y�Nx?��{iDb���ԯ��&�Ԫrm�j5q�,�Hb��B�X��ܑs��t3���
i��Z���v��.95��h���ÚĖP�oty4��K���#־�,�]WS�����&&3��!A_�m��������n�Y'U��Lbp��<�?�<�
�c��OAxě�=������U�{��~�7��V0׍��@Ɯո"�2�M�ӭ��ߩ���v+��n�
]�����h�������cLY}����6��15׾O�#F�zS�!`2�B�j_��"����"�2��`!�������hX�%69�u)�����`.U%{z�&�}�z�j=�����J���jWJq��P�m����ט�>&�g�=���V�������_��S���Io��o3�қ�hB�� JZbj��G��da)�gcvU�c?sW�Ƴ�@B��Q�]٬:�Ν����ɓ�x��%
��H'^��~&�<��������](g'���>���}�r�Բ���<O]���3-ݗJ�W�4��CU � �1i��A�K��#�nqr(�KL�$�k}�H5�7�Cٛ�f�~���Xo�����p��<�5�v�G'��_55	�e.RS�}�D�8�eIv �l�U�6e5�4������Z4z%�eDe����� k���7?�*A㖡u���
)��XlxVHYEB    3375     bb0߳����F$���Y� ��es�{	�CIVtH��iL-����Msd-�.�nA"R�w�5��>x�JͿ%�y�.gP��[F0c���4����ٷ�|��j��b,XzFL.����Qg�B�%�5�����G9����۸ԩ���m�~��X�׈��f|�̓v�䚨��5b`�`+[����ג����l;y��R��6!�y����2��
Yl�G�ڐ�8�_������x��LuFt��o��T=g�#K�|2_d��A�z���N�Qp���B�� �O`���`�Y#�*w����l��g[5��Y"�T��z���~�CN�8��Ci���-N����vY}�JIL��h~?}d�|�$z�r���{�s&�~�D��|�g���^AY��J���A�L������%jn���'(K����\�lZ��R�Q;����]�Q�~�8K�`��w*��ڰ��m�??����<��I�C%S}�JۉUˮ����s4��2qb��C���
�S���	:���\�\��*&m��B~�܀5F(�EI�>�i��^u�&�t�h�(� 2�W�Z$��� 7�7"Yn�e���WNέt�L��9�'�J�2땍"���O�?H���GF�����g,�z�Q�����6�#�,��n���_#&6L�"��Q*���g>S�3b]�v"��<�W�e߱���S�9ߍ�%��Bg-/o��J�!CH�A���*zGX��
d-F<�����G�F3.���������2�&�9<��{�ϊ�а(��z9����������?�B�Z.��?��jG�bW������ʠ����9�ّ���Z�N�E9�K��4R�Pa��p�^<�Y]�R?��׹�����iT;�oZ�1��I��{�����`��A���*^�������Y����ᭅ1}S�Ky�d�����e�n��i�k
��V���d��h�~�B��:�\��C���h�CˑY�Т��.���P�~�{7� ǵk!8�tA�X���o�Tw�A���e}�'��M�o���@���ǒl
Cb�?����	�_*��uI��=&BV��f�uv,Jn�?�����"�iE"�,@8ب��vQ�[�y2ٕ��,2��Z�-
3lT�F�c�%B��j>��V+ YD�ay4�$e����@�G�*�ͥ=�7��vk�l�SC��F����?53�ʝ����#�s�s��Yj�H�|���q�ӹ�`�M]u��o	���_�d�r���9�GH�)|����ց��<7cc�3�]��k��Y`��榣���k0������#2�Hu�f֥Qm��S��x�V:�Kǥ�L ����`·`�Pw[�ѽVo�-f��M5��t�P�G�V,B)�����x���+0:,0X6�O�!�L"�	�ET����7�ްH	�'���U���v8:��mc��A�p��%�l!I�Vxk�tޙU����8= �>�Y�yau:Ȧ ��bKz`m��x����QNz��$���5�d�OM=����B�Ϻ��_7�T�αX�*T�W�h�ѷ�.��zc����w�K��Oh��&���6�f�{,��z�)��Q�?U��������v��PW�6��%�K� �LԔ�8u�v��Ea�!&�2������ҧ�0%��/,�]Dh;Gq6�ߣL�;�ٚ�f=^��|B��6'���������K>��He<}��$�����C��#A�����������p	4���}�".��'�H�|���-��&`[D���������]�B�Y��u�+��AO�6��B� ���ӑ�*�RS2�����,��`�����9]���7����	�wTZ����'��%@�P���=���T�M,����Cy�h]�����M
���.�7�(�rH��9j,�׊1�U��y�;j�-㡾�)�@O��994���`��=.%J_WJ����t!�_b.���G������$��R A���o����L�a6��d��|�Hid�dg���1���:���9A	v�o�1�iڋc����8KG��:��8@�nz����?��>�,��D�ռR?>��O�3N�Ԩ�a%?8�.M���Jˆ��C/�0v��X�m~*��a��������Dq)�oI�mK"�Nn|�æ)
aYa��3�*��w�!��b��P)��Z��Q�ɽ��A��U�2�!����F�8�<��~�V��dq�Ɩa|r�d���ڮ��Q%݄n�x��:c4?�zw��`kW������_~��:��/k/b|���Xf��s&��҅�_��I3�X�\��O�p%H��AR�
����a.�z#$[J��͐Z����pp\�j��X�>�[����$@RO_����óQ��e����2bU��#"o�F�T���M�@�l$���`Fo�q������t�Omp�%�#��4P��޽ah���=�d� ԩb\>\3���������T��kiWW��.��u�Oaŉ�xt���]S���o@�1���z�@r|fL��sv�j' ]/�i��wqܾ���i�"W62���~��T���4�15J�,�ԡ���|�6�<_�r!E�;�$��&jK�η-s��Udy|N�`"a����"�u��C�-�фR/��*����^�Q�Lq�'��ً&𠥩!�&�����-�OUb�i)�d!�ZNn㜵�I}G��y��y'S���UY
�u���Jc���nx�<���l�����i���\|sOSiu�atE	Ӣ6K$*�|�7�a��E�����_�L��t���*w��B6fz������$����T�R�b;l��W����jƧ2��;��f�S�D�@^�1�S�������r���D��R)^�8��EPx���y�ɮ�FFa��D�L�8	jA��K�'X�� �����?囄���H���:�m�pv�Ǔ�d�X�:�Q���(&�]��?�P�78�	�����٭