XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��>�:b!.?/��f��o,IQ���[�3��'���HH.׽���a���e'�0%�0.r7�Rc���M���Ѱ{��#��e��֬���m]v����d�O��ʓ N�\��x�f_��2�C��'\���J�y[�Z�&�C�ǲ
�!���3g��B��]���8�Mۦ�f$Z_���U��YE�?�	�t��������{���ig�<�����oUTg��H�0ǹy	H�,x�M)�5q�{^(�S^�ʤaNe�n��G�c����ze"*���n(�Ӣ�o{�c��CuHd;i ��g��V���h2�jo�ϕNZ�nu��Tq���V��A�d��W�Ѥ��Z95�`��w�ɚ�ϡ�H��՟V��;3/�/�/4hQL�Fe���*^��߽a��L>-�mk��Ho�L�����N�J՚cm����4�K��4�W^W���^�G�jZ)�|�?	܁!�����
h���v��ֿ-^���	K�lw�yG��K���%�8_z�r�ٶ{��"�� w��<�B�	o�4���-�)��A^���-�#����E6�|�ڴS��jT(2��v���|�:̗*���l)��D��A���!�/tv+D�*H���%�r�p�.k�A�gըȁ�:��ו����>�"!��hz�;�B����8�Hyq�6��0�7MHh9�,�1�	1x����?�&�RI
|�Oʩ$��(#/|�9�k��� �=�n}�֤�M2&\XlxVHYEB    101a     450�����o��B��6':l{ħ��}��M�ڼ�h�'�� "L��+-&c��.��_��1k:OUd/_?a:V�.[��*�g�|��C�t�G0lpB�c1�X�,b~R7i�K�0]��9Q�0?&k������h�)�Wx4?^��l�~2�y��c;��yϵI����ㅊ��A�龩�5���$<��Y����+��G��Z�CB�olØFA[0�/W#Bb���?��7�F�N����ϛ��2L�]��J����?�߶��sK�!��1�����|�Y-��jd7Kg�q��$��37/P23tUR��҃U��f�_�X��I~U�1�A�y��]�s�.L�Y����˟:#=�����A����P�x�R������KE���M��x��p�(±M~�s�Ѱ��.y�@��[��KԦ�FH3Cw5k�-�� ���x��ԙ�}j5>�N�	e��^F�����w<V}��G���bꀗ�t�(�v��a!U�` ��'Pk�uj�-𚪳�4���; ֠뙨Ǩiߝ#� ��t[�٠B�&	��Η�ƋvR�,F���ᶷ���wn���D��Fo�|�����a�	�ô��'��Xp<<A�����:�W5��6��ıA�����Q�~�3�wWq��88��u^'&���#��9�!�D�]��g�=�B�\R'D.C�J���:�%��;�*A�`տ�xD�?D�E��4O�����o�z�Dj�z��rp��y�^P&bT��-�S�X��cr�(S��6S,��F*�Ч������owq��m�%�z���D��t8���ܭa P�$�� l|���둺� h-$��{y�iL9��+~��!{�ys�N�����D����(XF&�!#����ǸJfw�'�bwSG,<�#�+@�T����mKV���X�ۏn.�3g^HU^u�����s������0a�[��k~ܙa��YZ�~h$�ծ�YaMUUg�N/��X:��x.v��q��� ĸ��B+���\rG2�w�t���,����c�vb�H����u�mJp��_{I����8�D.&��)�����S8���cX