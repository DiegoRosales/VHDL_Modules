XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����Z 5a�Ŋik$�M/�',J�ʷ�PK��z���d������TS��� 勽71��*O��q�ي�q�8�^������B�h�pl�����m%���z����T�G,C�M�	2}$@i7ȍ��,�Ҭnݨ���*��&Ʉ\'L�Ȣr�C��&w�C����F ��J�0��r��Y�%��" ��'�)�NvV�vB:��P|����[c����t����Ғ�w���t\�@����#���!����$d�X�-ŲrK��Kt�EA��Ȁ5���-��ת:җG�\��Q͙�hA�r�9��>�#i-�(|�|����%bK�A,9 �����Ȣu,L��A|�����[�z�:YPM���ۃ�Ҿ��	%�u�)��S����[LD�����Il��0<�{��g AP��œ�W���,�\P�C9 2��3�?d0��pF��2��������0��""-y%_�`����Q�zd;�a�V�b�EHF]]��=��u.U&㍜���RΈ���40*@.~�坱�$o'����W�f�̳jS��@Z��n7���Vq���ݾx��zӚ
cݝ 8f!w�E��4{����h�D������*Ս���I���^�Q%2Fh��L'��i�� J��K �|��֨&��o�oI��TVD#�-�I��y�h{����P��X��2�_��lW�)Nej���P�Ū�_4�
�q4,fP�Q$�}�[��	�[��х�r{�6�j�{oXlxVHYEB    1264     780�T2b!#G}�8��
u*�uM/��Y���������>�r�@-�/7�{���� W=Ҝ#�����>x���h�Ch�2Mu��7f��@@��?2��?G�+�5�N����XL�`wb#�ȩD�Z�r�I�`��/�
�}T���@TRٯ�P�*�W��fށs�qw@X&vG���=���)"C�4����¿G�[�%��������f�u\�e� �����rA�*�ِ�l[�3mŧ��l�{.�J*���m��Տ�)Fw���z6�k�O�S�4�C�Na1)T�bc�v١Ҍf!�PV��%Ii�0(K�G��\�L;�s�|N��n�G�b���V=��*�'<R�@��%2�)�R-E�:�6g�����Oa����ny���۾�n�΅�6�O��{0QC���X./m��Nc*!h�ݬ{`���L�%k���H���h��P�W��BM��EO�A�x��Yq�j?㣰t�*?"�(P�7KN �e4��0��'�3g'�4���蕕SìI���/�-��^>��K�JEc,������.y#նۈ���.0���ƮIr�a��ʞ_���s/l��V6�:G�H����?�"���}��"]��8e{���!��9���;w:q.쭓w\�
���j0D^�]����t2���1N%O�A,�`�Kh���A�X�T��L9�Q�1 �rY�^�@I��n^Ͼ��2,o8����nh��2�YQz&i�+׆F�ݠg�&]���r����<��=�j�w+Wi�����H��~>(ֹ��M{���o]K�
�\��<����}��荆/Z1�vfx���~%9��i����۞
ؿ��������Ӷ��!�jx2B�c}|ٜGWy��Ts���UH��BV5|O;@��f���S�D.����n���۱��!	9�����ӄ�������^u�k>i�3A}A=Nn�(P����]��5s4�.�v)(�f�f`s�������Ŷ�����}2rp�^��K2�n�J�1fu�a�9=ι�n��5�4�f^���S�"b�������qi�nEb2Ɨ�K�-bE��(c�!g1v�@>�mZ����s����-n+�%usG�����]|Г��ϡ�O^��w��#_��,( �����#�4��~���|����x!�:����s`�VD�і9��Mo�����L@g琢����pq����V�3�<p5�+�a(j
e?=�"BԩE��f��\P����{���R�e�t�� �������BT��TeH�R�7��`�m������U.�}�����w�]T�0�j��5�6��q��`���;$���O+���G����IbZ�n��P�ly݆In�x��&�R�x4�D��^yR�<���3�TJ+3�&�/$T�b��>4��+4�$>�	�|���7���O���C˸Qw0����=}H�ld���fō��_�|OBK���d=��=��7s��6�,*L7�q�!�f���� �y��D���;^:��}�oj�I᎔�]����z�%�"�����.��ċ O<?���Kr�:Y�=�o�V%�R�"�G�Ӄ��@��jw�p�+����Pj��h9�9�Wi�[>U��]�)6�!�i#�C�\ e̃TQ&�@�t���`��Yt������pn���woV4'�#73Ic̈�I� F����ls�`���cv��i�~Q%$�M�V��?���ҿj�E��S��VB䜿�y1��uA^uv3G��f�lE�Q8X;�՘�����&2�G=]������B�aEƛ��f������a69���=�Ү����o�a�LS��54V6 {Y�z��Mev�����:~H�X�)��s_��i�iV�4��sd�