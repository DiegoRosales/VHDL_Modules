XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���-I�v���B_�C��g;��A@�~�0��Y	RL��W�t9�3v{��5!��j�~dk�~e�/}:,'��n�ڑ�iK�D�e��Ї��R�x��k�<Y�Q��'�Ғ��`f��t�n<5������-�=��K௥Fi	�Wŀ�!����2Q\��K<���{����=`f� �A^����j`�w���+Q_��q�j�U����o���b��#/�����D�w�NX�6�~{��D�F��L��:���Iϡ���æ�k���ڠ���gr��\H�Ro�Ђ��.�n�P���3Y#|�����s&���L��\�Ppr��bZ~��*�m���ӊ��7.��E��F�c/"�(���c�@H[�gv�O���.<I���2�'����2�K��>��w�B��o̜��G�KQ��OƏ1��@7���L`s�����A�]x�=��F�)�mk �_Hk�i� 6�	bKC�M��S	U�03��
�^0:)RN�0X�'/>e�B�S�Q�h43��)�R�΄��F�m]O�p�O�[���'��2tqR��i�ݍ���MAToKu/VD���ڸ���� �g�����#=�C��\�~���̷�	��z0d������L���q/�s���.l��o�.(�|�!�����BX�1��h���C��:+mn��"�l�0�D&oa�e��f>�@�%��Cb�q~	�tk�1t�DV��i�냥f!^����0�d�;�:ׇ���þ�c����G�G���WXlxVHYEB    fa00    30f0**8Z@#������+���g�1AA&)sĝ'm��d⿸�i�:�������;_T�C��5k�#�7�ܳ�26����Ń8Ml����u�s�^p��`�h;C��fῊ���mNT�2X�]Ch&`'���K��pW.|~��؞g��������F"�'T)A��R8����2l��?Y�1j�OX@��.�}P��8"ƥ��9a��`��Aw�J�~�� ���K�����^�ǆ����2/�S2��#r���^��>8>�.������1-$I�sg����#s}�o() %nI��H ������rK\��p�B�_X氥O���j;����L���]	
}c���-,O\n�~��ߺ1JO4����#�W��:l�Ϭ���������C'�d�+�Ī��_�yR�qy�/��f�=�}�Y�id� J.�Cg��)5W�WL�kQp\�֒R4-�B��l�a��S�����>���QN����9��i,zJ�x:�q+�!�Q2��pdc�B�vA�����	;����A��3����]�|�!��Ƕ�#�F�X7�P7�>YB�w�������OA���&o��(�f1p%��W��c���{� ���o�w��\��ȱv��(�t�i!czK	�[b��H���z��+9��P�d��Dy9��fx\hd��oT��{�W���m�7���~yu���h����l�|0��^���y�/�a����e��r�=�DuX+��tm����1��Ւ!M�C�]R�^ ���w�;���f�LD���v�Dv�t{���'���*y�ä̖_`P����b:@��y�ﾟ��.^�9����`��m�ɫh/l5��!������x~'�&�o�A��u���W�S��I?����3O�W#Ɱ7��N������%�6� S,�mf��A8��6��-+�`���%��H���N��N���'�c�Y��iaY��8�I,s�d��f�׀��Ѹ��S/|H`�5���4��
��Zk���^-�����R	��:5`ă����~[2�+تvT>i�����J�F�.�3pro�����Ew�R��M�d�;`v��᣻�XRO<�n+:��4E.��|�E[���i�p�����"����v�����<�~V2���mݩ1Sw�ZȭgG�)l���c�n6��%���ӕ�l�%�T�\��\oI�&OW�T:����0���0G_�T� 2�!��]���H��"����=�]g࣍�\�\������o�Wܦ��Ox9"��$�V��3d>)1�I�S�����Bx�~0	�S�G�Uc���[g���;���{#Χ��s���<����"6��le�{%]�qwg����C��4E�oPM��q�������mL:mK�;��:�����d=S��ƒ��3v���'�1"^�u��犏�QsiHqͰ�틬�i߷|!Q�7���J���.���G�ZA+�lX^^�I)���|�Ej ˗:��Z��QN�*�s�٩�!�6	ndʖ��VR��i ��ϋf�uT�"��^�&δ�^PPI�^�_�����#Y�N�����_Ih-�3S�� b>�m>�\bH�k���DL�da"�ISUU�ڕ�=��uqx�`4�9�{��tz����gt�������z�S:�YX�iyԙ��ׅ��@��'V�4N�;5*<�� k�A�gH���/�9F�2G`eC,A0mX��J�t��-�F��cB��Pϧ�]����,7|>��� 9	ސk�"׍��>���/�b�
����%����F�y|���oT��ZR�=)<;�����&zYx'R"�\�U�lx�3������KTd�L��-Rb�`��o]�u�l���_B3�N�W,�$�9�TvA6f���Ďޅ�D�f��H)Y�@��*�C1�����������R�x�r��>�6eF�g|E���/s�FH��>��x���&�u(��(�g,k���ji��<@\�̨_;�q3��6G!X�<=��6��T�M��[��cX2 �Zp~�ڴ�G�9�e*�� l��!�h�}���G��������B���q��~e�ز��:p=\�T7F�*K��?aph3#A�_�9�[	$)���gwډ["'�vym��N�c2y�~��Jw��y�P��N$�Xo*��%Du����I����Ǟ�g�=S�>�ڳ]�y��z��TI�Yz�j��n/1�ޥ���#I����m�"�#H�2�"Te�y^�%��В�-�,��4��5�]���.棓&A�hpmD�`�Fm1u��?Z��M���[�*6�A�">���!�C�J�&�
}�������ҋ��n �X���`\��B�N�c�|�߯�RJ�F��Ӱ,��L�9%U�A=%_���*���T|�7�S�)��K��c=���yP�������\O�SDGe��Â����u����8�x�j��
��~�qI��k�^�}�p8GK�fg�$
>k����!$�:���4�	��0*� �]u��uR��,��)��fb=PGḿ���B,ix�G����|��Juw��|(EaL�!�s�ߤ�E�o\�N"O���e�����������\8���ɯ��ʟ��i�Ih�kz�QԈk�,�R�sqK��t^�*Y�2��5���G����b\R<�,����-�c��Ok$��ڟNm�y,�]�4Z�0��X�d�8�8zN��n�����z)��E�n�C��*v�����,��Z���ҋN��z&n��H�⩄BxM
�� ➁D����y�}:C�o�;� P�
��mc\�b��*���-W���Ľ�ҢԦ�;l���b|��1b4��dXc��b�х���j�z�b=?N1A�K.���� +�%�:�o��W[�Ϲ$*��FO���۽��l�������d~�krh��r���}�{��]VuDs��@�oDJƃ�3`q[�7�#9�;T~+!����5�p&�
	8<J�3����C��Qa��CK[ڼ���{x,�-�iz��Wצ8���1ք86���&.���HvV��%q���?wPB#;��Z��0�����um$��MZ ,���j���W,E��w��c���2yo�������@�Jպ壒5ݽ� 8��3�)1H��A��;Gįs��Jd��ᶉ�gx��*��B���+b��I"�B����jJ��xq3�&]�a�֝��~hN^�v���������V��I@e�~��c�̳rީ�Ѹ^r���zF���M,�4�B	�?^IeFLG?�O�?�c�[�?)�}����Z�bG�2���V��hɆ/>���)�<�A�`B�슲�����I��L}ʟ�-!d�R���<z�5 �E�-��gPFm��w����m�h��@��K�2W"�PjY�z�D�y6�#i*�7��Q�pg'��/���s/r�����͉����Fw]����U�t	���^D|�3���5i��a96~5f3�p$ߚ�{:��J����M�0�����M�ԉ��?Q]���%��$�ݪ��s��	��7�ڀa3�G�fD� �eg_|��f�'~�0U5�k��j6C��{fK���km�<�|�]o]��\�X['O���Jb����[/��O���	M@+t��=�H=_�����e�c
℉�ҁ(3��S�_��t_|�'�*���F�<W܅�Z���kR^u�Wٝ�#�)��#_���Y��%~�B�`5�Le-_�eK�/�E�jW�55�@��s��m)-��'��F�����]1р3"���V0�b�g�@"���);`	0��x�=�,N��R$��0=l�F���NI�� ��r�3��Lkn6��}̵>�q���jmb�l�!�͘��;�M�u��L��w>��x���%L!��b%��,���y�Z.�bVG���<&(�t�	
�z�s�h0��Xk�� m��o� �&Y�I���և|�*z���[��;�8�t�������.і����t�U_o��T�]57�N�L����ְh%J��Sv���OM��VM"�|�[�\�mf�b$?|�����F�+�`����>�H����&��|�b�vq��Jy�]D�S�mh�
���i��N%lp �$L\���;ӝX�ØO�$��Oo\M�:�������;��lH�ת>��5��B1�ܺ��@�W2�`;c���T�WE1��r��$P:i`N��^=�|nTP�
�R}��B3�o8��K�"�E��d�o{�΍~
:��B^��N�N$u�~� 
�|4�2 �_H@�	�iH��U�Y�@��b��攈�΋�Ӗ9t���́���fz�S|��k��&���τKfC�BQG����f�R~Ni44�����e��@	�E���]zϠp\̉;7eWt�*3�FǤ!:flᭇ,�����ok]s�:޻�,�R��a�Se��$颊~v�
d��d��x���:��{b��Bӊ�*dt$~ۜ�t�=77:�k8�������P/J�]�x݃��?j�AO���Ll�8$3�ʃ���A	}(-񭬜زj8�uz�0���E��|�b�;4\�� i�������t��7+;8�ן�,���T~���>����u�}c����Z��>��ߊ����"S�.�9�ɥ���ѣ�'��nF�[e��d��L�#���K�hG��y꜆����4��r[3F��0Y{؋>�N��q�`
�݇���h�o��m����87'�H(	w��ylś�t6�h飄UÉT%��B�&����4�׵�����(~������]1���}v�&��C��(�j��j�2�"p����3�B����x�|���AZ�"��ũ���oJ�-���7Ym��z�͘;_�_j�O��k��-��B�vë���e�d凵�4!xJ/&���\�0���M(���1��i,�_�{��N��sժU�n�B��?�3��K<üauDVjZ�Ӓ�πoι�k���$U���"��,�Eޮ�],8@7 �� ����{�!*)�/�-��iESL�ڔ�0�$����>�%�g�8�ȍ{����c�vG�`�DD�T�1�
����3�O���2��f�O��L�|M�eIZ<�>P�i���k��e��$q�H�������j$%g$�ݍ��hW'��#7�(�U'MK���`��	��99:9��U I�y�hg����U���u�KF��� ���C�M�\��2��p�����H�j������xϟ�8�V��c٫�섖mje?:p)�:I��8���Jt,3I魤���3~�6�c�{�&^�I��8���ڎ#�IX�k ��G��2����;�q�Pِ�O�8��z�����f�8S��P: ������T�3����X�[ZW��=C�4�2?�lr�Q�H�������M��@�k���%V&��4Feޭ�M�Y.џ�h�x�l���>����Y����ݠ[�}ݒ�+H��B�p~k'픅r�i���З�AS�R(�5U{�&}�IS���������1��K��zLZ¦P]:3i'�Zb;�˿��*¯2�y�	h՞+V����\�c!��Zg�p��#�yp�M��șÕXOH�]$���yz�':�
࠾��8�<�@[����n�9t�-��-�+\�~\�b������Ɯ��c�� �,�t����kCk�|������z��Sc�zJ���Eљ�E���72Gw�C��
�]�#*)�t�&y%/-1~��a��em�a�%DK��+�'�H/�.�H�t�e�G������CS� Z+*O��OJ�<r���Ð�����Yǁ`��%w�ׅ��W2�#ݾ ��4��������SSѕ�������ol�	���Xk�Α���Gx�wc�Z��bˁ.	6�C�o�i&R%�H�7CH�Kw�Ǻ��1����_�R�%���Q-�ϛ��V�C�� �0�#K�B�4";J���0���Lj�t�f��<��x�* �U���Z
l�&UzΘ�o۾6\�S9�� �bN~R$�c�[��s<�f\BTE��-�/a�G����O��,6Y��6�o�v	��*�����u��,c��P���l��[�㍟�`���XE4U�4����ë{ѕ,(�
7�$�a�|�S��3����[
O���wr��a;�1>���E�Å�$Z�Ũ����(N7�G4�G�d�������`���3��U2�Y�EV�_xÄ��	s�G�%��γM�1�����jv��R�p=�"��+jrL�qꔺ�С�A�
yk�O
�iHg��q��K@RC$M�u�Qy�3�s.��d��������1��v�J����}�3��N w�o��~���	�c�ޙ���Q@��ƾ)G���T^/#f,=�
�y��Ҧ�� ~�D_�\nk��H�Kʫ��|���ǭ�m��?��-���8?��l��B>�.ZZqh� >�&K3��s��a�ϿW�f�w����u�״�Y!�8B4�FH�*آ�w��kS_��A���{� �f�[�Wθ�:�P�m��|63"��}���C�ױ$/�N���&8�.��6
D�$K;��k}H�~�=wN����n4>#S��Á��wvd��D�E�8��5x�T.͕�U�O奷~�Ȟ�1`��QZ�8��$uV�"�q��J�z.2��Fx��y5��rܫN�S?��e[*�{��jǐ�˅ �j���A�5�S� ]�%�ޟ�:w���Y��=�J��U����#)-����I�튶R��Qt�R�[�԰��|<z�:k(���밟�S��5Y��$�n����9���P:�1���(�/�W.�	=jz:�t�M��Ο��`K� 8��!�}/kt�l[�!+�UTcה��tp��N���(#W����L���\V�D��&��T.m��4�� �̋�?`�ރ*��s�?
�9���8P�P����^��@���Fރ<�S:B�{�W���EX�4���b�K��=7]�#�az�f��Mz����ՕG���s������6�N]��s�Z�)T9;�귷C@�� ���[��by�2@�7��8i�UqHղeu`m�:{��Y���y�䶌�cR/,�5�U��,���b��%m=������ݛ�T�	�o�P��X���
��˚ה���5FA����p�<�D���\TI����}�Y��Sj����������4�B�����"Uњc�H;�O̸�8�U�꡼G�7���P��G�v�Q���m	�	 ���vRGϱ�V�t��u�������G����b�e�\M"\?O��kpOޡ�&Y���]8���YkrOZWm���$�xh�_�;����������L��g>�
��l_aA��e�����o�%0���+���SOz����"Ǘq�]`�M���a�9����Rhxm̈/���Z/T����:N��B��u��zT6�74p�j�y�.�$��Iv���iޞ2�(3 ��u[��s' E��C�E5����"�j�8]��p	ŀ��{�\NqF"]uOz�y��W<�J��h�"ࣱ�klU�R�ç7c����5�dϝ�~��B��.�ۧ��:_���m^��ŨB�RRw]��(����^�^�g�:������3�Q�]�3��k�\۵	b1_���s�U�)����O��`�����CyU���H,E޼Y[�X9ib��7�ޓu�L����3R��������|����X���,��z՜����앃��0*�ۚ]�q�K���9�Z8X0��\\�9��v�؅N��z:+��5^�����hU��I�
��*/�ؿk�/����m�?��kU��uC�1G�&����-6?P��ꑱJ���=[�?b�Gy����s�[�*��Wk;��v����(ଟ���#��ƫ>�/�d@F�� Hq-)*�q/�CCfiv?[��}Y����.�i�dY �= +������w��@�5�X�~�8>(�?�)�[_Ia��#�QNBu]��hETb|  ��݉<�{_V������j�G��;�ǯ��qTe���]����+��r��vz��+'ͽ��9@C#k�$N��Y�}�SNΖ�ve�)H���y�a�����+���AѩK#������@��;G9�K�ơ�ot6w{��l`"t��,��j	�y�ķ	��ߧ�� q��4ڭ~���+�V��j0��/����׼����< 6�N�}���/0T�t��K�ҷ~��&�k�Y2���F� h�{�So�>���eaE�����e�.���h��TFNfq'^�!�؈�i߆ɊG� |��;�+O_�@���>'�"Q��*��激�3����ڞa�C+�D#��N-g��s����/s$�jb�Э��='�P�BQa	c���B��8y�1�'^)y����aX
m�Uq�Zq���'�񫚉`���m! w@�̜��~6" ���bA��Ƥ
���B���A1��O�W#��D�7~���<i}���ڦȽ���#��u���E6f��,_��\�C�#+�xߜwBJ``LY;�,`s˗m��}����!��$���ޑ��TN ��`�����H1t"+8H��H0$���hzt�h���S�e�������ar^.�!�B�a��pu�*��Nř�e������=٥0&*�|ed�W�w>���M"#�/�<�2�=ۤ%�����Y�`$͗�X����) ๗b�C������FmF�׹�)l���oT�"#�n6C�j�s-Q�
�dbH�l�w�`Y$wR��9������/ẌV��V�.7�s�|� �Mm5h�K�p���-;ُ>��'zu:�\:7#�jo�zH?X��t����>�0�N&��5��/���R(I����e]�k��9=��z�ce�p���bGy���8��o$Ǳ��x-���)o�d �@,�҄]��u49��Q։�9�̆j�
� LqN�FL�^��ً�}��Z�:����j�f��c38��5�����L^f�6s����Z-��xtΨ���[�a�h��G)~>�;"��ȱ��_� �4C����8)�}���O��e�U��_T�ws���0��Z����LC5ļ;C�Ō��k���P�����h4f�>�hwXD:NMh帅)rCG��Vu'$"�='v�gF3�]4.�Ns����0;�v�	��b����]�V���ۥ�Ȱ��"Q�MT��_�rF�r�٘��"3-����v��iް�6L�+���cH�����L3Ԝ0ٮ���	{��\V�v����H:�X�6u�ܾbf����ܟ'R�S��$�=�F���J�M'[��W��|(pf�٪���[����x�\/A�sߡ�]-4�6������,j�9�Vp��Rx+]��3��f�n���J�y�-��#�r�E|�`X�I"��LP�������nO���e'�J�^T���$LK2�`d(����1��s��i�O�i,Y���_F{��K�>'e�=���:�8"������{��_Ơ8B�$��tc�jB���ay��Ԩ��K����.]|O4�=����EI�/Â���#7�	�]�qj�Wʏ\�S��q��˱l6�ly0S�=�!zI¾���~3�Na�{�rZ{S�5�hG[�z궶���y�%�Wr���� �`Χ�0��y���<�R��Z���sS�+h1��Yʂ�6�D⻌�����)w��S�)��˻��� .i�����Ӕ��BO� ch��	:�sL{C)KŞ���Nn����)�o��u-t�~�"Vy��~��AU�H�4�S��
W>�#a��G��?j��Z/�To��M�Ï5@ݬ`��%�3.K�F��j랴�ŭ�z���F*�Q�s�>�B�D�˕D���
�֭�b
��ڊ �ƚ)z�f��'����ms������xc+x���������*$J���O�¥�u�<"�����IWA<7���B���[M<Gͷm�%�p���F	���d�?K�#0%�E�MyAɎ%��}�&���ɨ1�z��'�V��UQP�����O�]�pP�ti%SE�L��d�(�������Xc�
��~�N����`A�H�hlf9�.��=�!>L�)5���U{::���MΚ��L+�wA⧰b/o��,��}ޞ#9+�����{Ȩ�=�z�ut����V�ax��+l�Zi�q��Y�%߿g��i3�
I����8����Ú;h���u����a-�g�'v�m��nNνZܱK�P�6�Ӹx�N���9� ��|��r�;�������8�W�Dȋ~~�kL�:O{�ƭ~e��[P3�}',p��|��/*�t��H�#���Y�����U �{T�o�R�3���
zļ'?D��g������D��]���W���y�ge�N�L���+�����p7�Gl��J��i��e�D�����):'bMa3
�s3o1�!�x
�	��\<-�u��5=����ρ�Ygd�B�I���Al��w�zGa���z��a�z���cY�z��Bk������+�hɨ�Q�J��R�� �����(�9SW�4��z�����Ԃ��������E�����2��? �8@��
��w`�@��^, �Caǧ:�!�rj�Mܲť2�{C�u�FD�Ut�Wwɛ�.�apr�L��?��v��I�P�ea�����_���y�<c܏ ���2A�Pb�|�P�&$��,Ŷ`0��|��E��������W��4��puo��-�;���`��K��9��DQ�B���k��_$;ߚz&���dQGӅtA�^o�	�W�#�vMOhd 4�9�PB-m���'w�1��Fܻ́k��F������}�%��"�q3�&l-��PS#5j|�N�w�ū�bⅪ��m�s��G_W���g�ᷳ�ʏr�&�[��>�-7�{#��
9���-�ew�ߛ8�RjxxOg��Vx��Z��.o_Z��;�-��չT'�c��;�c`�2X�c���d˝k;���oJ��J�|�U���9�V��P��n_ݤ���C��:9�R�W�Z
Tp�L�����@8�+,4�WNo��&v���P�� ��}U1VlR�"����XE�آ��l��u����OB<x<���⡎����ο�����+�_ۂ�J���Y2#w���GS+�A.R��Pq���A�?���/�`�����s����L I����w�ss�2�-9OhP;�3�i�P�$'�Vɇ]����R5��w�{��D��(��X�u�qu~�ra0@`"Ɍ|���ة��{�A�U�\��Y�KV"2|T��cm_!���b������Դ�b���7�o��ա�H��_�;e!�A3�P^Du��������Q)��x�����������F�{r�e�ߖ�'Ab�0#��d�@?�Y����f�/Qo�-�A��6�e�S�~Ĩ�}e�����c�ľ�r��s�wPC�_��2y�����,/�|:6"�߾�S�%/:G㵟RF�������J�`������"��O�2��)o������)��Y?�� ���Z�_��iO������0"���Z�D�Og�<!��]�_��[�+��������#cRRCo��Ψ"�m�P��W�ϱ�"�:�R1<n�c9)y���Yݗ�A:K�t{�d±&V���X<�-�M���^�l���z�k�*��riq�1���O�ݬ���V�c�%�)����CW|�ӏ���ci���Ek��Ԭ����c�B���4� �ft�.n���Eʋ��f�(!��49�+/�J�.M�iW����+��[#��C,�N�q#��&^� 7Zf ^��H1��Bg$�-Z����	����b���	��E8/�[��x�Ǻ�����^��L�����ذ��W�@'JR���\GHJ�S2�w*���l�T_5B�k�W/�r��Ȥ���KƝ*FX���J�̅z1Mc�Nβn�x�ͨ��������n�@@�q��F�X�
���>�^Ӕ|���v���@Eh-�&VL`9^;��|tzbhv۵P6�K�R��O������IS�/J�H|y����b���)H�U�I2�6/���ƥ7"��a�H�r��_�,r�#O���g�nAH�������(��>ȅ�WOf���|��U�x0���'ࢊm�T%���w����Q,��̴}�9�v�8�� (�y�ɤ�Y%�=��3vHPl%��AXlxVHYEB    ab24    1af0ȏ��+:49�B��1���Dɓ���<�@���Uv �v��qe.�?�0���8_7:�1�'���z^������o5 � �ք3HZ%������c��h��N\�"�@�RX$��������I����S�4��	՘��%��{�baca`���4�+(;�Ki�Ia@�!\������{)9�����u�ǂ�af<�
ԧTw�*���NUͼB5�"�A-d�����g}���w���,F�-<So� /��$�H9��֐��ѩ?Utq��c�S��:$j�~F���+�JV���<���i�tNl��c�ɡ��
K�8���|$�Y���k@ь5jWS�!���>d/�٣�����?��r;�4L���r�Jy�R�F����$ߤu�[\q��T���3욅��3/N�L��7����ap䙉+B�rB��[�_`�}/8%ޗ�*n ����XGO,:{�����D�c��y��A��J��dƁb��K�Q�ɫ��]�L�*����X�_?@:Eן:��۟>yøx����K)�H��E�;�z�k�����<^Bk��5 ���9�4;`|�V�!��^�W��%IuT�9����E
��o�V9МA��ᙜ'e�}���eh^V����>�����t/�2��T8
����Z,Z`�h�܎q�jyϙ�R�,�,gR۠H����p`�ԌPL����K��|�,d��	ix�d�����J�Tt[��7<���}A�B�j�M�*eI�ғ*aEשS2�L�Y��r�&�'*��^���-(�i���W�0�3�lf�A�?U5�k���)��LӨ�����_E6ɬ����Ӟ��U�Ӎ_����R�-,��Z��/�}2���|#�Pg�8��ڱ�6mʾ�pJB�O��2��yo�G��_8�"}����4�u9\�^ǮT|IӪ\3/�f��n����_fH_�(�I`Ӎ����	����N��`W���� <=!���D&rvD�&c�����Q�D �ɸ�{#ǚ֢ u�÷ꛄ�$����́����Ǘ4_'���.�!�"��Y��H��x
-϶��k�K�ϻD�CY8�y|p��u�ZǪ�A��K�
��m(�E�) ��TA%O߂���������c՘G\B�������l���F��j=���=�w�M��- s4�7�4��{�(�rm��V����Y,)�j�~�7���o�j'�Y+'�[����C����什�g~^��m+����G�p�SB���4K���3:8d̶^��čXǼ��!�����d��vo=y�B����l�r�?��g��U� 9#��S0�xbe�ov�����%�����q��T̝u�	��eh4��
p�[��o�-R������g+.սs�����%��2��`I(��J�԰���ÿ����Ϗ�/K�U�����]n�N�x��_�g2�n�	U���1T�������!�x�L�;��8�B�jN�2<$�ӋN��Kx� D�#:�Q�m�ʜ����DW ���s��"i�jCº@���P��-k"'�8��9C�#]�����G�}�M6��N)A߳{�9I���@
���Ľ��=�̛�/�[3+Sp:ج�eCP�����:A: \#��3C�:zu��I?Y����o��n�W�@�/�����k��ʗ 3mF�zӡ�t)E��
i�:?�TH���!
hJ���o��3�ڗ����4gE�-u�VɻiyB��ꣿ������i,ש�-�����S-�y.5���U�g�8����W�ROj�ٞ2"ٚ��ɾڴ��N�H�*�����l6�1xj�/\aV�]Mޑ�p�.f6�1�����:�m�\�y�ɪt������mGh��zМ�ʾ�՟�ԙbt�wS7õ�}����'f?�#/;��L�ன 3 =�����G���hbp�0P�n���쎷)��Y���+u5&[3���ӗ1߄�y�gQ�0��k���oU�vS�}�S��1�55Z=qNJଈH��3��Z��G(�޵���cP!)i�
=\�B�3�ik(�҉bTy@��U��������6n㿔;����Tp1��Z���^f��z҉�-[��m�|}��z���-FN�����8�X �=܃C/[F���f��p�4���]00�bz����+Qٶ���F��(�_�/�Ϣ�����~C,�!N�����7����m\�KFQ��L���h�׉���T�RBEv�	�C����!�?w[Q���(H�}��:>��6�Y}�S�9�U�m}�l,��b�!9[�K����F� �Ց7���/�'ȗ}����.]f�a�!�k �6�wҹ	v��f��6�IP�BM��	���urq^^\��z�6h�׊[��{�:̥%z�j(V������
��>~��18x�� +'p*c|&�Y���3Uk�w�軲I���s�0ҟo��'u_��4m"Lf� �~e2�ʔ��x����x���xpԼ�S�2�>��q �Jf�[���J�Cw�3�DW9~�1�W��R�1��eA�0�%���S���D
����s�v�C�/2�����A�h�?0����o:$���
dQ�jfsEK|4�&dN�7\�L(1i�&�F�hZ�uD[T$!���p[�����g�(rW;�)��.ǔ=5�Xj࿨G���%A�+U��}��CH6�_�ʑQ�箦��9��-��~P�D; f�9L1��/�2��t &%1.:uthЦ�,Zɋ�$X��a�c�V�i�!	�+&����fz��d�g��t��~~�S�`D'��d�ۭ�41��5�j�-^v �|ϝ<Y�H�*�`.b������0�~4�vm[F�ַ�B=tE鬃#�`e<��HL����I��d[k��=pp��Ȇ2��G=]s�R+����#3تӖ�����uC�F�^���܌����/:^�(8�v�%L�;W�Խ��J�ޱ�mr��1I���1N�����؟6٩�4.��5@V֛�\ϰ=���Y��qB�����S9?Y��{4��{>dR��21��20ϙ8��TX"�M������2s#/$=���jEţ�G<c�[�7̐)�a��Bm�<*C,�g��j�6l0j�����;F'��{�F<��]�з����
��`u���#	m�p! ���U �ԥ�M$�/����g�2�][ H����pm�-�>Bt�zPc���w=+��;�w�mTS{H�5�T�|S�F��|b���1���{��]���/Ĉ���c,�[5�����ܨM����k�� ��0�O\���9(�{}W�o<�'<���3r	L�1��Y"F�������i�/����3� On�
�#�qS��5�'�t�q�7Ve�s��h�K�P���� m�}<6�Q��#�b�ǗԢ<�ۼ��Ҽ�S���b�0�\�Z��p ��j3�/��Ac*~�� o�E�u�Nr�V{s���'/H�;�A���"�U��v�'^�X$;M.h�w��$2st	�!i��|�Ǣ�g\"���2C~��V���3 CJ��韗��Pe����u�d�r�NK�_}?"X�V��`��	�e�ND�3��5.jjt��Lx�N3�M+>k����=���4~�p���������(����c.���8C1=�ё�\�"����0f�5pU�#��e6��v~��9H�(g�wCQM�y�f�* ���³M��F�>��G ����"��D��w��t��)�.Uae���*X��
���47�_BSƈW��
^z�6�,7��7�Y9��$7`@�E�����+`�}uYI��#fTjY�%�I����Nj��WzE�-6�������WF�W$��ރ�}���-eEʆ����x�=9?bݿ	-��?Wݮ���R��M/��L��31�������o�	$�����^�q��M�����+�/
S%0��A'�6���fB��Y�(T=��2�[���JGm?Od���~���C�������&L����W�b�����ڡ �F��`�c��ӚH����I���2���.F}|��y&B檬2(�g�:�������))�;d��:��������x�(a�ݳ�Ƀz��*�x��V<g핱��A���7�ݕ���iS���P��� ��W;��_临�8:"~��j��:{<�,��"��Cv��9��Hf��J/�pU+���"�� j,�)�|-Suu�ʡ�;��I���5x0~����
�?��#��:�LC��P��_%��-PWpAZ��!���>�ج�僉�s���SJ���\t���p^��Vq�Z��r�Rk��d����3���p�~IJ�o�`l��:R�]O�w��/�-E�b���ũ�9���-��=�Jd�I,�H�p��")�A1��#��(�9��K���-V�#����~�6_C��o�� �j�� ��F�m1���1�hb���;�d�,S�A�l�� ����xQ8�l�U�%�k!S,��2`^���s������P���bs9��H�� ��@����XEf�=�pym��3
9|���x'���[zI���`b�0�s�	Pxм}��+�Q��ff-�߿��~��NA#|��J
R��0��hۣ	-�i����:��q�1�M%��^5��&��f�ٺ,�����ݥN�GÒ����
�h�=?��c {��)��ae>����S�� Ւ&� �B�D2��e�a#�n�wr.g���B)�P��:;�"��d&�Kz��@���Q�<�!�<oP�m��K�g|��gvpx��LMH��t2��7ֺ��<P�(�^�`|m:�e�91�g����W>�B#�N 1�8��hda t��m���=>w��IGh��e��~x�v���g�1<�Nص�v�Ꮀ;�,|S~��	�n.n�Lۣ�ć��[܎���iX���v|FY-hn�H��a4�f�'@�*zQx�p��?����LSM�d��Zs��(4�C�Wi0[�%�K8���sJo�;�HVa��AVR��oܗ���0�PU�l��z�z��q@^�W��0���G$�1�����E�
�+G�c"���fRpGS����\=�8kf!q6��<xf2���%���i�ĝ����%��UE�<���	_d������ 4��>���
���^*m�wZzԇ��K�{ ��j>g��h.fY�k��;�W�V��Z�#8����uE����2�����%�	���u�Ƙ6����T�!@�S�����t�X�/,��ty!�����m �9�uQ�tX�d��.	�z����7e 5;�ѱ]��A-�U������2���W�,���ּ=$��Gj���z�^�HB�|9��.��[�ȉw�����U���*��ֳ�0\���{_����<% G=Y�-Cutu���ҵ+�T��
P��ˆ
H�-���*R�_�j�K��>�	�IDw��o�D��>D��b(J�h��#E�rr����*E���$�{Ѥ+&�o����ZH�M�m�qx�grlt;���Tv�V�zi�rڜJ�n2G|9��o���T�~���|;pg�8����#�|6�Y�r9:���:�z�=5��#��I�=����h��܀½3���}�H88�|�5��wʸ�;+�Cf{9Ι�6�,�
��(�����x�NuG5`���� ��Jg)�"�9���*�O�B�b?e����T{��Z��)7�	Mb�Y��s	���i.`q	Ũ)�P�e'��ch]>4I�M�ÝK��=��[�]��������.P�`|) "��qyV�`�xw\����v�JH]�ݯϬ3#���k9��+e.S�tjɥ��n� ����4�y�"��#��;h�&�1#�j��CiÄ���4%rDx��ԩ�r��	�`�(�6�W⏕bq}����Z/ +�k�t�G�۞(��MQf?�%�Zg�7=����umKc���0�i�Z�[o���`���.����dǄ��:���������y��2��">B6cL[�i�=K[��BU\����sCč_���rm��mU�T�B��J�ޓD�0'�
1f�h�S�h�HȽN�ǚ���e��ǼK�ֆ0l���D����U3Ư���5��M�W�Y�W" ��5J��XS�*�K�X�ؽ�|�5��~?�DI�H��ɂ�KD��3�����7ۗĸXC*8�N��ۨ�;uƠ�P?���ub���D pѤ�X_�qݏ��ŨWy! ���W��Q��ǀ�lFiFŉ�ʹ.��H�r�/e�z� &��H͆����e�y����/���j6AD�=�{��^� ���HmAV���<�#ޭ�<v�,Vy�~�Yo�5o&UER�����������Ŀ���Rk����F� ��O��I�*'H�=��_����*���Ե�M��-3t�(��c������`�[�����o)�z���M+ˌY�*G;����@�B߹o2�y˹�=�L�=`�'����m�M	�:���H��+, �� �U�Y�aZ�|�Y��`CF`�oZs~����� ��)~� �6銥n�T"��u��4Y��:���H�����B�,�&ry/�f���S�$�9  �3��<���� �@ ��tkF��^����ڹ;�q�i��N�-o��JVG=w�[�buźӭ�?��2v>�ݑ8<�h?
&����Lf�Y?H��\�Dc>S��c���v�*�S鶤�
u��N����^�Fn�>IR�����YI��M��ߩ�l[]����|0#La���Vܱ?\���i�4N�L��8��.�(���C��m��3Ċ��