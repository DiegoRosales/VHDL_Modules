XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�����s��/&�x�۽Q�<�M��:Ð]6����,	i�ȵ�Q��,I�F��P��=T�/���]�b���iIU? rn�QPm�M9�ȉ~�;~�&��%!q�)�P#�v>�?u�_f���	y�n��V+4r>uD�n���T"����-��\��>�"GB�b�>�k
6 s�{�%څڟ�Nqc4`��<p��Q&��|����p�y	�4R�k9ה��S_�����E'e
�������+&\dA�DX���65�s:0���5ŀ��3��M���������+�p�)lB���������m����*D�3�j��&>� �3]0���2�n;¹,��{�������ao���</�I��yf��đ97�ၻڬe=�����+�@=��d�KA���cq.*�T��E �`Y-��lஏa���+^u �~�xb���;E/��Q�r	� C�����ԏ�0^���9�x��eRc��o3�<W��}�`Ѱ{I��5 ��6|/�b<��U"����:k\�kLE��H7�8��Pت�@��5(w�"@�i�8Ц�7|����w�)��>���չȄ��I�ag4�l;G�&<���e��0�-ۥ��
��|7r�zA��C,�z����ӳ��k`��x�f_��D)�V
�.~�	�nk������(���~Q�^`ڦ���^�������^�>@��?��ʁ$bYD�\BN��]��8C,|8�+7��8��瀬��+ӭ�ۀ��嶜�XlxVHYEB    fa00    29c0�D��/�ۇ��6���8ƈSUR/�^R�5A�S���V���JQc���BT!���z�=`D�����J�߀����A����Mh7�y� ��`��(;����������.�o�%�SW�	���7+ƊdL�oK��8���&,��g���1��+.~jl����Щ�f����g�tg��Hr�TY���ʔ�����8��L��#���fF��3d�߼�>�WSC��5�_������:j{�H�w���eJ��TU�*NU������F��Wss���<���x�5�,���(�m���E�ewi�P�=��yQg���#N{�����:����\�LMvA�~�f"�ᙲx��U�oG�ǥ.\J*ȿ������#��$��h�h[��#�*7�"܈���7tw�Mp���'Tm�,�Ӫ6V7�*h	�m����D��J�Sy��^�[��Aاo����2<[[n8=�O� ���_�O�T�p��z	�:���l��qkq)L;;�/���n_�Gۂ�e~Ȑ�w�/��)��O�����_
~lY�,p0��Y�>z�#�y�'��o�e%�,ԙaƅm�fa�]X�kW��HZH�L���L�L�Ŵ�R����q4���Z�ᔐl,}e�w��!k����lE�3�u��*�c$��#�����H`u�D4{��gS�S`����`�=�ܾ�U�G߰6�⒆ �>���k�h���v� ���q�'��!r�8��8,��R��yn�!�,�.�b�9+���ߢ^�^�k�D��D���{]�g���&G�G��0u��ݿ��4�]/���ڈ`�l��P�#���bmL��ޒ����
Rm��2ɯ-d���_�Bp��(<�"sk���-�ȗe��ű{9R��>�b��S���%n�P9RH���i0��CS߄@��������<��J���N����<3D
�d�Nj���#�pN��%=<��ɭ�p9K�+��2I�e��k�C�V�\)�O�� 0B��k Ve�(��������$�4��NNWxI�f*#�f~�!�tp�T���;]�����6L}�W���@4.��@h�q�b�&+�W�܏�E�&o@��>�1V�6@�t�L����8�#��.�F�}�s�񥐖냶������c�G/e����oCd���z��0�������t,.�*���)�M�ǽ�/��m�)�+���=�`���%cF�#;Xo��{Y�[�b%i���y�ޟ��
H*?Y']�%-�Y�~Դz6�0;G��7R?�"��3qs0P�����t+W�N�u j�iq�",96�ja��~W�d`im�6�,���B���Ɯ:���6(�����I���G"td�ށ�./���/���3C�"�����
=�;��]g�Yb�{��t�J�86O�CFD�a�X*�s=��׍HǷh�@��SqU�i)G=��_�P���T�T���8L����Ird<�W��jX�R?����~�(��Yq��j��Q@Oct�Q[����G�0��MX�j�X6�OU���D����<w"������	ԍO�ak�[�`��Dư��]�jLx�d��qmM�l� �˙l<(=��8O�c	!�=e����� ����W�$ P�:�f�����k���]#D���&�\.�H,֧�7(D�M�����0[
,	I����N2���`ck�F��R��i��*�`��b��qWk�B=�;%媴C721�#+�:�\�8���B��a��7�`I/�4���*[�p�
���u+�Y*����CJu!����'�[�)V��u��P �J)ym���s�]�O9���`=��_�/��)Y���[���jF�ǐ�VwEI:� ���qQ���	ڐ���T]���;+$R���c݂�B��V��sv�m�oϠUQK�?����b+B�#�'��oH�}1�gR?Ё�nQ�P�!�GJ!`�3Ӕ��y�?� mEQ�0-4-�=�pb���@b�l6)�X��=�2n�]E�;�!��)
��	�����1{��2�����^}Yc�B༯EX���؏8!f��#�it�i�V��N�l�V�L�/�3��ih"�[z�����A��B�#g�� �d��wӔ�A@H�^{}�8��_UoťVZ��b�� ��ae>�Ȅӷ������4*G�-%f'Y���{\q��S\@�f��\��'BH }S-����O-�;�����43�=<)k���>�����+��5@.=��C��7� hk�D�bu�*��.�%� �s�d/"y��Cw�Q��'v6q<׆JOcY�璱�K
�{��0P:)���p�"2#�yT��U�S��r���'���$5�|����؉5�ʪD�t����4G1/�$�Cl��R�JJ����E���(-[�z��5��Q��|j��-/�=*`�����J̈�خw����WE6^lt��������SS3~�# �K�	���E,�yIO ��w� T���Rg�其��6� O����ɖ3~hn�&�zˮ�YS�[D��_�L��JHpS׷ʶ�u���!���)Uݕ�;C%�7�ߺ��מ�##��[�
:���xQ'�g�PP��QY��� �V��+�s��^��E���I���f��}�P6S�g�����j���x�����U��^������4�8��T�#pp%�tCW�j��p��)�IŔ�2��%4�V��&zs_�V�[bJ���b�ZT^A�Α.�I2H6���'�loj���b�+�~��Ќ��B����i����Iݧ;�������qt�G���y���=��.�1`�)��,�K!Q�De���Q1�|�D)%R�~z�w�P��j�0��\��_ˢM��)�ۯ�[���Т��X9�꡷,f�_�t����J��P��eR�wt�pTe�E�gq
����0���V�岗/�#El�x0�g'���,rTC��o{������������,J�-c�7R9�
��:� !v��.j����:y�Р�!0�ޮ�Æ�d�5g���X���L��n��B�ݞfVB��TU�(ƌ�
�߾�6��d�8��#FA/ܴ�=�T��}%KΚ�uk���I<�:���Ĵ�hCMp�9�n����־�=�q��&��Pv�����Z>�mȟf�5��D:�[F�%a�+���g'�5�|� I���4���[~t᜖��x_�TLAu)97�~�x�"Qu;
�ON��{�~� � �/P�9c�'������h���5�W�J�j�����Q�uZ��Zu���3�dO�3������4���F-Żs6��϶���̛<����լ=e��.w+�l���)F��c�9�ʵ5RV!7؁pO���d��+Y���OL'�ijߙ�����f��Hr�A$��ao�9H�y�T+��O���b�
 �c����� ?;a��'��.Վ�֞
	y���e��]4��rmv�F��`��9�>�p��ڼ�X��,V���$�����T�����]tp�?��6�.�����M�юa�����.40oa�Z�vܿ���rv�T����ҿ:�%�aS ��aF �Ѩs^�������5��[�R�XE<#m��ؘ@�?��C����-����6�S&�s��3�[л*J�L��x;�+m3�hS�\I�:�é?�k�u�~ӽ���K0S <5é�R�S7XS�኶�p�/���(�)0Ic
��utK�\���a�y���c-9�l�屟QNZ�|�.���ɅH�W8B�DVK��d�Jڒ�Cz��`�,�ݯ����[��a�s-ȋw}��-���=���x�툩&�p�슸�P�#��4f�X۩a��7�ץe�j�Q�PCR0�y����Ÿ��>�Eρ���M�
����L�X��oS���1��"��JPe�qZ ���:��k���4����K��uu����ȩ��޳��o���N�n$��m�&�޲�Y0��c�b�X�� �u��Mj��j�! Yc�j�n�!����`�����Zې��}0�?>�Y�sG�}|��*}Q�v�Z �W�䴯[T�(�8"��,���N�B<z,o��0V�]��L]�P�X�'N�������I��yG� Q����Y$�LNQ"!���^�k(��3=п�q_,��������6C$��i���ñn��J∰\�m�*�TX�
t�kQ9ެ��:�,��m�|���H�*�LE��lU��C���z&�p�u��>oZByq�.������Ԃ�޶��7�4=�=��@���ؾI�����'�*Ce�p��q!e#=��cP�A�	%״�]W���͛r�=�k M�>����({�+Z�ZG��"�
.��E��ih`?ڤ��}�-=��y	;{@$Pp�,J�:$GsC���3�1J�����hO���O�ʼ8�g2��6��k|�N�AĠ�U:<�y
Q�Z;o��ܟc �X{�x,�M�z�ND>�| ��sv*���#H��4}��"4�g{���T�<�DT����5 ��(�����,���vȂNE��PlD�9��6��M�����Yy6֐��Ίx�8h[�����=/�t�ލZ�Y����~j�������:b�´'����6{>�䴹��!đ��y�V�!"�V��ı�������ֈ��C	2�B�{מ�Jt�w����ĵW[:Wa٬A��9;
ܔhH_L�zo��Q���������\���Kꔔ�!�/�o��B���ZS�h�q�d��a����ބ��XU�խ��.xk3#�f]�9��x� G�JmnH�c&8'k1�Z3TbX�4�����C�'��v�i�J�@n��Y�-"�Sס�?Oگ��(՚!*�$zD:"��ND�>W�q�^��g4��l֮��yK��{>>V�P�vf��~���ܬ	��U5�~��t|]d�Q4��A(w⒥�NOp�",IXA�����Hi9�?:��x☴]���j��f	w����1gf�r;:4����9��,2S��w��K1�6^z �1*��<VMn���{��!���.�W}�I�xƛ�r։�N�� `�9GQv2XPU�G�i���ŞM�i'���[F�{�E��6)v@?#o��,'4B��mۛ��l�|3��uY^H�]���U���iS����ܧXw�X�e��Qs�/�I<>Pw��xڷK����y]�ݤ�_X�����[�	/�5���ٮ�P��ڟP�Y�M2+��Vs�����u���v��2`2�n&-Fp�˜���:}u��?�k��k���s�P�{��,��c ����jZ�.�-����� ��f��	�?2Rg��3S�7<q��T�F�'����o�º�淬��-�'���I���0�S���_�rH6��e1�MNM3�t�*��j[��T�k�j���y��4��E8�ы}�R���v�5ƌ���k�!򍖲@��MC���u�*?�Jq���A�T�j5��Ӕ��DyI7NƝ_H�$Q�sƀ~k� y9��[��t�8�l��X`Fv=a�?���U�[ƺ�Z��-h������8�@��g��D�f̷i��I\�{��X�+�/���=�6}j����kr7Q�$5�s#q6�
�8g�*�@A|Cf�� C#��"r��?�����&�ϭ����nl��<��5����
�����!G���t��°>kV9��/�4ՙ*�+��x�j��a��U���S׮���Z)�"�4�\��g/�K�-�Q���2�QC'�wR�(�sه-����i�zb��'J�B.�˥��$�No�X���J޵�Uc%�A  ���Ֆl��+UI��b�i#NVp�h�MF(9jw!����ƞ���q�8t���|̣#2�ˣ���?�@
�'`p��� ���^(���}��H M����F�_�\�sA!)@Ŵ�o���MK� ��ӈ-��c���F |���r����;��n�$���j�G�j��9V�`^���{Q�)�$學g�ʙ^*6�a(
I(�I ȔI���l�ṣ�n�J?" mR�y�@H�Ǣ�B�ܶ }Cɣqǖ1q�������2|��	D�^���
���r� `�ǵ�䕓���}*�ż&��FRE.�����i�+�,��<��E��>o�>��`���mކ#�����w�#�U1m�6E�}�!�7�٫y�l��R|����
��>Z�E��b��*�çJ8H��6j���������X_K剜��;]��ϔ�L2�(B	(�\̌;�_X��$�O-� �I0�hC� �v�������R��j���V���`J�!���#:)�r$�j�}*���#m�n!��G�'a��(@e\'��_��p,��Jjz��WUF��K���na4��&e�yV0s�B�^�����	�2��髗�+y�����c�gtd��%e��qN��FZs���L�����/^\�;�V��Ћ���&��v�=���N��{,@���s����D�QsGo_�&�c�G��$��B�Bҵ&���/�*���b��� �_7z�:����I�!�~XY`aF5l�u�4g��t��xm��E���+q���l��Ɛ�-�K4ה�?��="41D�$���g�4��:� �?_ʆ$g��&Տ��m.Kh�*��o�	�;bıfn�֪0I�I.�2�������l��l��Id¸���z1��HD?���kS#>�+�6m��<��0�cs�Jo�x��jTª�[��#z%R������b�v C�_z_���y�Rɼ�ي�9�*Վޮ��x�~Թ�������x"f�Ծ!��}'nq4�b�[�N�J���ge���P�G�g�G��w��޲���N�u���	�f��6Nƕ&}��~O�޺��X�;x�u���jLAp�9Af,)�RW��Aͱ@�4�|(c��(��s{tf&z �r�fa��jo����0`���a֎t�>�C[:5S�єWJu��������f�($��n/7q�v���\g�6���vJ,-�/�I7�U�^N'�}-!�B	�W�VX�g�Y@�6 ��C;d�GH�+�c�Y-A���6�t	\���� +D�\�P�}�裕̟�/�vR�aɊҵh
���@8�)xe(G_�hv���7���Km9�~*����	5��}E	z���<.�'�:���)�2G/Mv�nf��;w���|�VP)�qPV9TJϮ�}��]}jބ������S�"%	���ǩ��p�b���I�*S�C<.��W��+-�� ��n���M���K^�����ERK����c�S�l�КMx�8��H�b��T���bb2$@��ˮ# �~�#��� "�G+�U[�1���ŋfݯ�u�m�m�ܼq�K���G<|���g�I�:�gY��M�Y����X����i��zw�UG�� sL7�#xR"eg�����Q����9V�o	�BQ6tT�\�.\����Ȕ��턉��^8��\)]��7)�̱	�]=� a4Mm��C(�M�{X�|!BĪ�-�$���h�����Nzzb��l���E_�Όַ�t�{d��k��D�ʆ�|��!P�&�߹b�\��� ��'=�l��)���♢�e���`��l��-�����tT�)�9ӽ}��Ȫ����|�ì#�O�2Yd�F��YX��(�R� �^�ϻ��đ�)ilW��Yd�r/�#�U��Jn���=u{�m�l�o�����?�IH�vH����P6e�I��<�_�Ī/,��%He�;�,�W|c�.���-�p�M�}N��c�N��_ ~o�qO����10͝uiޔ�e�B��V������ߝ+�.����~o�%�mV��g�|By�װ�j��n��X�A\r�<�1ףߍ*�b�D�H.��hʼؕ���t���c=���g�7�1�^G�]<�xtEVX������NS�JJrAj�z�����n��}`��QT`٘�V�§kܵ��ny�jH�.��w�v���~1��[ywN�u+�p�?���Z���FQ�
ZC�t��UZ����~9�G�dd!���9ۥ��AG�+C0
��^�G�:EE�5΄I� [����3�7_��֖�+,�s�w�ݢ���vl7a�P�������x|k��xg�����ӗ��g{�S��&1Fq���� ��p�d�@z�]��`�[����Fĥ��l���(p"[����)�%�˝ '|��ۖ!�b�W�C5�n���4�M�O��B4-x��]���Q�=s*�f�NfYU [�TE��c"�6��w�K&`G'�g�cQp�D ��e�z�p�n1?�Ϗ_שp���O��h�����$W�g�V��^�Ʃ��=�/��;C�0l�ڛ����=�+j��C˸v;xH���;��]�*a��Z�U��8YvQ���e��"+���2�Q�0��J������eq��JSL!4' 5���:j��o������x����r��v< ڻӊy���	���.%u�<��+��.��0(��憰w�'E�Cl�H��U��%��ە$�2mB��V{1�F������g�<}aC��Ю}P��}O���e>Ј�N_���Q�S_ds�5����ՠ�q=�����7�x��
�ȨE�z�?ܰ��3U:* 1zq�����������dU+�d���{�s�LNǻ��PV(���;�eJ�%U\?8y�����j�Q��J� n���3z~:J��V)	܍(b�IH�Wg3A�f�{�"�>�
�伲:�~���`���y��b�'��)����Bc��h�k�Q׊�M��DI��|����]>�Ω�����\z'9��%`�K�Լ�NÞ�o�s������ɔk��Ӽ�ڈl o��RE.�C��_LN��R�6���&@ ^2wJ5@7_CQ+c�˼��u�+�:n�Nz��o���9h�3�ȧI�n!L��T�o�M�O���w�i�C_K��`�7�Y���?�GO������Ӓj�3�40�<b��f_���e�0*T�e��(�`A�Ø	#�g`
QZ��9�� ��A�� �����(�& �;-Y�&��L���B)Vh5$"���v�d'|Z)��:`�ϛC����bn$�@ &z�C��V���\�緣ާ�"�nZ'���OT�̏w������ ��v����}&F�;����cAng?�֘\˅K9�ty-_�(���/"� �<!Nk�o�}�¦��A��V*LKW��w���x7��@�T9�K	c4�pb8�.��O~M�X�7IDr+�ayk1_� t�%�h�A�� ��W��oM�B��)���o��I�y�y���̷*���-bZc �V��!i%��dCK�(��URmF6f4���ʭľ]9po EB��tIdg$�J?���7\H�E9m{.E�P�+@~���R�|�����(m2c9ì�8�+!�	l��4wU�xx��N-t"'+!̈����c�]�&�M�m ����s��'}���m�f��`e���w^o��N�p��y-x��O7 �U��\\<癙���D�~X@٘�$�uWa�OofR�e��bģ����N%��]yh� G��k�"+ �RvzK��G4Hا�FhU�XN>r�r�|�hM�#�8]�eE�v)N����Sk��.qG#MqD�)m�n�~���6�p�艆m�L�ڈ�M�?�0�C-���7
�K��K���_"�j9�b�g�b������9R�wȪL>^7�� }|k=���
E���fg��)�/���"�ф�C�a�� �|@�x����[7�i���͑<N!Ͻ&�����r�P��#>_�T�i<Y>X�,��I�"�U�	��P�Cr��Tυl�G �v��v5�}�W�zb�N=����!�̭��R��"�8����9Px"~%�i(���ն�����jBf�����n�j{��"�"k`֞��O��'ڟ�ǒ �1
�N�K�@|5�П���M��9�F����E���	�R��E-�b�~���	w���@"k۾Q�ঐI�Mz���>�9���'byth.�z���5���h��¹��G� j�3���m�\Z�\h�[��sZS�B�C�gЋw�h�ک�j�y���}��i�~w�tL�8��(6�� �]�g�W�Eq��7�o>u�V�+��5�p���2G��,ˊ/֬���ސ�s��8�¦�U ��[^X6�Hǿ��[�]A#K�Wx���z��Y�`��W���f����':��>bQ��̩a���I�O[:|����V"���@�9g��`rخz%gٽ�2����Ϗ� ����v��Mz�9ĳ���U�ʥ}F�v����eC�:������|�Y[�@g��2r �U������ć�r�m�m�*Z&.�8~�5w����n�J��p8R��&#jq[x��iK�E�zq#�S��?���-�F��N��lHR�	e��,�Áa�z@�~ֹ#QxR�������)�߂[���9h'XlxVHYEB    3507     970���`]_���F[`�$\�8声/MD��ݴ]3�x-�?��c�P\��|u��N��S���~}j���t��,���%�
B��M-`�����#@#�U.��I};�Vy�Z�Xĵ�vy�Zv������R}5=�v4J���Ġa� �JwӃ�������>=�0� �9m�)p�w<-op�״���� 5��)q�6�-5�V��s7=��szS�|��:�{���D�=D��r��G����73lPh1:�2����L:���+�Y4��#B(����Qo�Qbo�Ua�A�6�,@�6=	�ekgG ���"�X-$H2C��	SM
d�ͳ/	QJH�0�s#зV������(І�zn�4���ٖ ; &n'&��9/X�_~�X�����3���4��8���W�.��D8�-n��XB�r/�!��H�u�(ea5 1'��t�d��O��]��f��>�j;*l�ה��e�+� \S�X�ʝj�(�ZcO,��gJ��^��g�a�Z5zUu%��l+v���<>]��t������>�jGew\<��J����o��!�<�qS����k�����N��)^]�2�j�}�.�T�����b�f]���q�r@p�Xʏ��r�oG�w��@Q��8"_�J��/�R�Ǎ�;��	/XΆ�~��w�/]�8�O��\5.~Tw>��Ds��G2b�s�I�2�\��w�s�'����Ğ���/ﬠu��[��3X3�Fx���Xv�h��RgGX�0 \�m��!R!��&�T %l�#����Q��`0�`�3a��JOGBؔT����`�}�:���+_�J9u�l�@��,�ӴsGEhchB7��U]�#���̀3)��;��Bm{ �d��D�qmiRy[6Iz#����Ը�zwpQt�,#�hՒ��ËG�׶���?)�1���`b���99W~d�J���I[�.Rn����눧�1i���R���ߞL|O�nG�c���%Ԇ$V�E�犣�Ru��lî��� ��|^���h�����=W�F������拇쯙 �-�k�+}m���T�da�,��e�P��*�>�{�%_�u�g��\��1S��f�	o�I�k�į���!l���a<:U�Q�Q�!/7R�����N���k�u�Vwj��a������[�K�ȣ�}���4���M�n�]餜�4�[_<R�������=*���"�@����{j&�hˣc��0�ɻy!pr�L����uuc�G��fF�?;���vեTݡ���6�7��jIc��ZeZ���&~�`���]�E�:`�]r 1�m~4Sp���.�R׸�`��T��K���\��Q��hxβB|W������8nI�E�X�����`N����C�2��vK��h�(��w��T()��Ky��o ��Cp̫��(��Ff�ѻ���E�7��}�A�`�Ĉ��ռ�{�t�w�,��"���&h���픛���Uf���E��q%�j������	�/x�{��^':�w�a��/�X���Z|�y�O$�{2^��^嫚(�Q�[Y�?!��#7�7�v�o5	݆m���z�ʾ����GB-N>	�Jd��N��
�gp85G�C�%kJ'������v�b��xy�ԅ���@\b% ,*
v�������J���+J�r�>��
���>:��.�����$�����D���&��� ms���}��=5~3��_�8��V�_ �C;���X��$C·<Z��k��&rr��9Z6sv.�},6%���S8�"���I%p�}k�G�)��ey���{%%\�hS�!7�I��:ee�aI���=�q�s@(n�*�}� ���}Y*{�4iу_���z�c�K۳a�s̭���f��i�?�<tq"�ը�=>Q�����@���?�Wh~��W��'�_���6rǫ_��&?���h�S�Dz	{�k� k���ob'(%%ۃ!L~s�e�S;?�&�����xS����K��l�i��Ƭ47��2�e���Íu�8�P�4$�ǜCMK5�D�Ǎ�{�N���DNӭ���"�>�A��d�*��`kIe��(�X�fhIHh*���{�f�l&7b�ϩ��i6W�b��s��/�&�-]�#0�h�����<pR��$P��i���ԊD�S͞a��b�&�~�/��7 a-���=t�y#�r\�^Z�@�4r��݀��/�l��w�a�^2B�O<]m�WJ<^����0Ӽ��N��/��*��`9�~���L��F�f8��A��ɷ����\=�|ߊe	�/lS_`��Q��l٥��oj�����=R�
�ބ���d��`�zN�I�u�@��
���C