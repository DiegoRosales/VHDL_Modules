XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��ezE�g�%Y�J�m�i����&�M�F�>�ij��'2�K��9�M�"��N��W�>���51��m�J,�^��F|ܹ��==P:��M��j��G�e�c�~��	�S�P%���ɔ���~�;�� ������F��;QB��;H�+�=ݲ����,�,���u��1([�����݂-��e�� ��1c���ٺ���K\���gN�'��2�u�p�΂e�ـ!w�7�e"O�M�A�4̼�m('v+� 0��Z.O�O���c�\79����0��x�{�`���Gy�:�@#dD�)��<�Y�o�X`�u���_���<1�bL�cX�P��?{�>h�ZkjY��!G��7��|�I��H��K�+�d:�n9�@[��q�Q��.����􈦛�T#�>��*�g`>g��,kȽ���)%����zZrRƁ��,�b[�&�2}1��3�-u�,L#x�?E��t=?2K��ˤdz]���
pd�x1�J��iƔ>����s������GX���l0�lek��.�)�e�^�W�Z�⭛p� ��N��~�"QTn�A����Bt)��v-)��Q��6��߀��.����<x3Ne9}�ٕ��+5��}��~lX��,������kx�-n_u�N1��X��Æ����&�*$�~��>�.��;��Kj
�Vb輎��9�rMam_�!�\%�Y�k��&�s��f�	��"�����z���c���ʡ��tqJ��ж�)XlxVHYEB    2252     b70rZ�ί��M��&�.GzU 2^$��t��@�^�0gK�ۜ!h����0�m��F�q�%���Q^��S �p�0@�{Q�y�I<ZBAl2C�n�C$� �]�r;}�b��Ť�_��7�U�I��)���Y,�����(�sF
�i����� ���F`���F�[Oz�;I���G����pP�q����MӇ%Kx9%=�M��J໒Ӹ���ل���'�'`�&-X:�	&�f���*?���Xt;U��w�J=݈��S���Fiv�t�6���o�2�͂Ycx��& N�M�~��8B#�"�w�����B�<@�H� ty�����~���" s�3�J��r��u�4�;v@�jK_*���IL��+�����Fe����\��N��nWM__\)_/Ns�P3���f'Vʵ��x�%����,����DS��Ņ?M��N��y_a"�&�g>�,�������%4p 1<��mu�7VX�	YN�L\�@�>3��dSh��K�"����&\Uc]Kp֖9r���-u@��G<���`XoXL�f)N�N:�K���R����h�h
�-��i��/���A%��@���kL8��f�8�.fd���K�ޚ����pƗ��|�����"���Q����n��?�A�gp���#�ma�s{��"������O�26��)
4Ju�����8m)��a��(���-	Q>f.����Kq6N��@����Y�KX��(UŒ	7&�2 ���H��m����P�o8����������6>{F����n�®dD�]�4栖�v�Q�a�6Et���w��'�jQ����J	���
������㠈�h+�p��
�9[�gѰw�^�y��^ܩ�w�k��Խ�P�o�z���{R[�r�N�������;5�
����ݼ)��L6�Q� �2�ǆ#���7�<aU6�ͧ�A�O��]���=��0o�$�h�|�#��-Qd�/�K<	�@(p��aapp8���D;Mn�H�^q{�I�X���{������ha13�ݟ�����F&&+�wHR��o�S��b=���/�Vt��%2Q*������.y�`����_i`� *&��+ܜA4x�C��1��^�L��e��� �	�T����Z���q����5>g�r��Ix�%)cC����{�O��Md���-���4[A�[�X��P��Y8Q�1���v='���T�e|�>��c��4v�'�M�R�[��Ʊ4�+��+xb`�p$�{�9b���W&"R|1�h�9\,��H\�e�S撄(�J{�(����ڄ>_��c <}ox��69�dQX��_9[��iy�)�z@��.&G]l�9嬐�Q��t�0�k��t\��U �?�콧$SM��ğ���M����r��Qt,rhW�Ky���;Q����! ������!���!�^t,�w���[:T��ƴLŖ���ӹ��\�t�>���sZ�2-,U~��x�Sfѱ�CH�Ϥhu�r<�H��u��"����[�����jN�*�%O��B� ���>�k�Ȉ9H�{�E�p��e�Pd���ű���i9�F��H$"��G�\���?We�NjBY�q^�M��`Z�D��HO켾$��9�X#yJ��޼=��b�< �r�F �������Dt��+�C]v9����lO���G�a^���&`��֬�o�A̧!��	���=A4,%���/*Þ���%�.t�:�=�1�Sc�c�l i�R���6��������>P`,%ْ]��8�^ܹ]M�
�@�'�k�39x�� ���NY��$v$�ځD�:7܅jwd��Os:Y,8�n˂(�ώ��	Qz-���nF~Uw:�i3��A�������Jê���K4��i���eW�c_�]�v	-m�'@���;�Coo��N���reUƷ}�6$���ʍ΋�0=��JM��=�g�ȅ�אP��ٶ�%H#���3
����R=MO��/������d{�����wF���Fv\"�g����.�Y��|ٵ�I��{]�|�F�1�	�F�*E����Ǐ���t�r:�����N��*<����$r{<i�Ԩ���u).���cRC������-4�`�����/A�^S`Ԃt����\u;���x��A����~�VbO��������T3Wp���k��s�j��C�yUj0K�g̾��,�:�����*Iy�\+�R���W�1�<�U_sG��5,���y��ýx�ݍ^��%=�3�e�+��Գ(I�,6�f�K&����r9�DU����9��.���BM��UB�KFU��z�W&��� ��������p�wz���5D ���m�~
�/�ԇ�VԈ�[�ӣE� ��'�ay,ƈ��180��������l\�J��!����i����b���U4A�+���a�|~��c s�,�����N��ai���B�͡1O�Lʗ�4 ���3#�'�����(�]���u�W�NR�"n)�y�4{�d��K��7������ǜy>阸��9phd�#���� &��U�L�i��g׾�C���X9��*@�,�~|��?tg���fU{8�[5�B��Y.F/�EW�l���}��#�W�s��M��{�ǳ����#���0L��l���n����Hq������&@��~*�~ ���g�׮���a'�6C��[�Τs�k�H���p���~�#�2i�,�R��y}=D����4a�ws�H�ǭ�%�Π�r�sƈd�
��u�	-�X'�",�mN!�ˠ��͔�r�B���-b8gU��	���;ߢ��=�R�]�+a������grlLI������n;q��$��*oȆ~SDk.