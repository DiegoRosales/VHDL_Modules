XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��S)Cwa�N�2YA�QH1i�+�&�rw�����t�2�"�'��b;wa^�ŏ��a�@6��$�������܌lbq(�#��E	���� @J�S��]R-X�MW�(-"X���{�o�3<����q-�BKv �M�7�jܠ �&<�hy�Z����*����Z��.��n�c9G��X�ł���2�.gNh$7�Y���������*'! ���Y_���y�2��?/���A{�TFB_�RU��R��d���oԛ�SÆ*��+�QǢ���]���6���N�l���)*�X�ʘRGMb�|�fd��6Q�!>�������	�O������_5�Cj���\AO���e��-����4��S�7�b�:�)�r�XH�g0*%���O]��i�Ҫ���9��Ï�:�~��̬�4�z/� ��+��.���63u�K�d����c��<�z+ڛC{(W��B|��WҌ��f�ho��9]����%D�#�T��h�"(iF�΂��Т�4ԟK\$XV?Ƞ펶����`��a(!��P�����<	�o��O�}�FE'�J�х�~�r�"�KĀ�Y��m�ѥ���
H_�DPŮ�,&
ߌ�ɬi�^pF[��*��n����e9ǎ�a�0Jf��8�������9�Ρuz�p 3>�;'p�
�7�$jHV\bV��źv����~ȩ7��O=.��,�{
�m_k�G 1��?!��d1�j�G�b[�1��k���KFXlxVHYEB    e5f2    2ba0N��ȃawj�$KGt���ƈ���ح@��;�M��e�~��
�D��e������xv�#�p�s��ӼՀv��o9�Q���yv��8��T�[(q��˙����u�5f����Qf��S��+�t�EK<h�F���*�,Ȉ|�����@G۾�t���:��<C�I�o-{�@ZZ@���a=_���@jM���}{L�J:�Z��y^��2S�D�8nA%
q2f$�Ԫ�n����Ѫ�&	��m->��cv�X�ɿG� �)cm�1ߖ��j��4 \�����ZV;��!����
¦f=�܍D�@��SB�6�Q���n�odAN�#��~๙�0d� ˧�|��`-�'�[�a�FV��59�T�����$��-�>��[���"3�2�qL	�)�^�6�e1�}a�����d�Q��6����{�pYF���,"�,#E�v�u.Zt�Z�f�M�������C�}�Pdt��h�xS���\���ݿ�Zu������&0uO�.��_�;���/Ղ����t�Mw������6M!�2��B/�.��Ǎ~��<)�u�a _u+�AO^RĬ?&rС|?�����g6s��^Xr���A3��aR�j���S�%5�ꫤpu|�k$���t�ėڪ�1<'J
1��H�U�����/�]8�{c~�Pb��ѫ�d�G�+�����ǜP�3�jijI$����L�i���� ��I���^��j*k���jg�ۈ��O���վ��9",�Fv�(�.�vG�|�A�97Lf�Jo (��~Y'T�?�Q�n�?o��#�O3����n�	v�Ȯz|�ni�aJ��W6�U<��C�vw�VJ"(/~�B?+u���ZM|_|�#��+����Z��e���e�Ng<�j�Y	�Q�?	��i��+�|㑓�	]�g���3�]��8}v��!�Q�	~�E
��1�.�B���ku7�(���z 	c'%>�b���%<�ǯVϸ��}n���\/E����u��f�A�F�+�E�5��� ������=�������A�_��ťq�r}�"�	_B@���zo�[-�1�jC��:��4�O�����w���=�����LG=����0$?f�'����"M?%�s���L��knP��	��A�������Г$����K1�gA�3|�4�$�ZԯS�r��R��$��嚓ǰ\>1���=��h��ɲ�G�p ���ؠ�
�I��ʕFg�����9j�%N�&v<9`�������U��푒��o$$;���ɍ�O� ]�-��5��4� �D���lv8�1J�^V{��s+c`0��P��%�����P������ ��X|!���r-)P�'t>T�N�4̵�C�^�<#!MT���J�sS�x��\$���굲^a�T(/�v�3iIc��A~d�H�z��#@hY�{I|G�`�ب�%�`ڟ�R�7���K�#��5"/,���@��������<>sn2_��I��o'ͣ�B��fK'ryM�Zi�/-�:WU=�"��Y��UF϶O����>bQ�v���MェKd��4�=3����@:�E#��Mg��M��F>�O�\=��<����cS�E�$������T��7q�t���H��DA��1�P����&� iڟ0A ���єH��s���Ș�Koz�dH8J2�Ë :���0�M�f�
VEf����8:'�-嬮�O�f�r�$�X�xP��p��)��ހB i������)x��)�*	0�x�f�E��#��^Y���6����'��h�@�k2�����^��ǹ��{��o��lT՟E�g�M
��N��!��q���ǟ�C��XtEOm�{�* �N���(:A����(�C���D�(]z��KR����P~י�42|Rd��8����LٍWce���Dߗnt��~Μ���`Zf���{��I���W�S��lX�����ok����˾� E�` tJ��:���]��!�%<ZB�O{�2��0tC�#��*t���A?@ѡ�*���>3���nX3r)@WK@-W�-Z�#�,��x	8Ʒ��ȩI{*�V�����H��sUQ�h�I~����7o�dNqB+��2�l��J!��cX���(Fc}^҇^'?]o�%�㗷D|��|�w�s��H���ɮ��F�OVɼ�n��M��]UÉ<m�b����Yf")R�u	�-U_+�27�g�H3rzo�*���|�*��1��?�m�9\Bm�5�[��F��Qzػ��W�%>�.Q��m!�����W�8P:�ߑ��"��_����c���Gv %���2��;h¥/
�����j�K��`�/k��΃}�`�v�����m��C�ϟ����Q��$�V�� �� ��؟���c��[-���_r�;s����S���[����*��63����U�ҵ�Ċ��N �nHx�.�*��2�U�w�3��xp燝�}Z�eGTp�'�8���(�M��.v#}&�B(���VpYݥ�,�Ru@��Y�U�:����>�U]&�D���J�B6�[}8�_�F����o��.7�a�o7mQ	v�H���U�)C�ɀ����WN|�2�q��~ad����L^j�����	HR�a+Hԩ���s�{���w,��!Z�+x3+ܜ�0����+vA���0=q��(}^}6���t�L�&q��m�^��2��Z��6��b2!�37#�3�Z�%����?�c�D8�����t���º��Kx^����n����w����JǓF'E�<kc��������>�9�Ӡ{h����T-pdtG�,���A�̔	Oq�3/�A7&�8$�ِ|�tؽ�������zM+ �S�+"�4���3�E��o���Y���K��[��uCɒ��eDZV4	��=ߪ��g�oA���V��C� 6��ϧ�ĉPJ����?�����e��*j��b�I��h�o��C����2HS;���.�9�C\F�!!z�����|R�ώN�o�i�>���2���`u�R�"��$�<̀}=_�u�^=d?�t���@�\6��+ʨ��$���	��	�����piOߖN�W\�P��񲀍��[�1��b����Q�{��L{�@Q{��`��Zc�e�RN�b���:K� ��&�>ڮL߅D�-�����:�^�Yި���ݓ����Tg���5� {ݻ�ZF)�i�p`
�F�"+)}6���*'�L�n���>V"���	f	g���T����O/xp�_�>�9tM��p ��U�D,�p,�)�bn٬ةvA����^�����5���	����]keR�~�*p��0�-�<�K�y�<��[�L�������E�����v�bAb<p��*k���,��8b�������������I.)���b� ��[%�8��Ѩ�V����$���S(Q�� 4K=�H�F�m&y�y5�A�!c�
�#;�ݺ/��GO����՞pk
��]a!d��\��m#-�Û
?sJ�乚"Rh�#�Y��ʾ����iW�p\�x����L:Ys5��3��R�;�	���C�����x�{:n��貅r����`߆���˕�i��t5��u���
͇&�.O�~r�kU[���ӛ��C.p}�+䧬�t�_n��K��������W?̗�f���Y��$EV�GI���o&��J��&6��c��e/X�̶�����2�6c�9�چ!�y�Ǧ�K��3�Ľ�7�y�,p`Tn�f�H���Z�Å���~����7�e�M�C�r��բ����C���g��b��F�x����@�Xx�� l/PF8yP����C�GB�D'،��d��>ĩ���|.�����P���t�A �I6��D�l��f��^�G ���P:Ym����
�������C��`_$^��O�FG��"�5�X��o?s�Vp��C����kxDt��~eV)n@E�,Ӯ茷�
����ˍ�2HHwY����C�f��u7���**$�w�!�8�K����8�o��M�v2'���clN�)�W��[�)	J���E�a+��_�5�9���j�u�P*�vWy�MK�Fְ��
g�(.��*��/R�S5�ԖTн�mA4ԗ��r�2�{`�ݿ����۷��j{ȥ�J�>�@���؎���2�;�_Nm����3�f��M�$QMU�hV�y;�]m�R���k 5���nS>�7L�S��L��M�<l0J��g�=�������#��0��/���&����{�.�T�n�$��;k���wŏ�,X"�.��R���/8�	�@��{nVo�u��=?.�)`��"�H��jB���ڀm�3��. ��<�qDY$��|��>4�(n�~+k��eu�aQX(V��V5L�^�)�1�(�����;���g�r�{�5�BY�wZ�Jh<M�{ʲ�X��-e��X ���j�/���Q�3�F�m�Z�@;�c�(g��f���o��}� ��fݸп���*��wG�O��ޤO�I!<+�M~X�~M��9d�g)5ӷ��p\��I�;3<��a� �!#T �Me�慁��ĵ��;s�1��hAw)�@[f�w��0A85g%a�VeU�PwH��#Sx(2q�4�	Fy L[d���G���H<�ۻ?��)$��0��x�}V�ۮ�n5(#��:�"Q@!a=�����C,�{R��*M̦8��N�b�e�'�v�Y�| ����#b�_������+h���8V�v@\,�K��Cɰs�W���Qd�L�� ̓��n� t�,GϺ_I��I�e~Pm֋�\ਤy�L����	v�����A�����%�咠��B�kD��{Ɗ�ޅ�R���	G,.Pl�i&5/ع)>�j3��#~���*{g��<�顓*A��m�f:����{2�sYGk�75�)Q��Z�QL��m�!�類e2r�-��+)x�2�=���5�3�MF�h�{C<�j���u'qg9�h�i�,�O'r��lq���0@�C�@U5v}֥�tG���0x���z�̨o��bU�ƶ��Ι��	z`��+N�Fx��nO4�C�k�������q7n�UN�;�ZM7bܤ��VJ̜���G���)A�$]�E�-&(㣘�#:�`�q�������#~񫐄8~�+����]͝h��q��5��w�^��#��� ��pS����S��,ec����/�V�C#�G� V��\)د�9�v8�ٽ���v�'����*�g�֓<:����qr1%a��9RD^K�
i��q�/=���w7p�S�V��O&I=[B]"��f(ՌP�$)C�}hXǼRuF� E��eϒ����q�u���F¸q�ޮ����Q�����~{�=u-� ��{ju���9�@���_�M�+�w�?�SC�v�Iȍ��evM�I���W���^�ց��9\`�v��U�+ҙ@ҕf^�2���^�蒳%��a~=����9;��	����"�IR���I>~!b����$��z�4�p�lܘy��2�[�q�^ͺ�@:$�3�+��6�~�
/K��éXR/h06|�l���}n;*d��C��e7�6LȎ_���`�2&V!��8��P@=ש�#�^��SV哂'�#ڃ���D��a:��Ԩ!,i�1�r|%�����!��Rd�{X��G�6P�{���H)�8Y���w�_Ĉ-���[{O�4أ	th&���V%�"9���)h���fa�'c
�K����R�^�q#�)\Z��p��)�$�4����kHU��R8P��qc��� ��fy���gַ�VT�w�8���Q;����%-��}�����&(�)A��KrDj���u�槃����!=L��Gh�'���7'���4`ؐU��/J�� ���=���� �� '+v�A�en��n�lN�e0z���W���	��=-�d=ZEb��5��n�rz]H�B;�/I��/��YH�\��'V���ɶ��G�'�u)g=���5������w��ٛ�؍{�i���^���Q��P�p�Q.�ԝh���%�Up�#��w	@$�{_����}y���I�����ˉί0������Q5�5<��AHv��@3�	��?��684�3��}{�EaƏ�+�0- ��F��t�S�mdL�@��muz6Id7,���b ��7=���� �2�1�y�.�U������P��jxR�� )=���5�G��/-��`V%O.+u���*��'�1��Ժ�7�VhfO�� �����>B���?�_>�EX�e�"r�BS�B�JטW&%fÞ�:�G��RUAe�����xmw���b�0�h|р���!�?�h����4B��{0�e��t����"�JV9��خ׳�ݲ���_��v��kTՅ�1<,)��2V�q�o��	�Nk�f,{��6m��_Q�0�w����ޅ;� �:����;���QD�S�W�T
�DE��ۇ��NKש���������6����h�|��%I�3@�$Q��"+�[=ou�:��~:>F�gS�����!	2��s0�2*KGbl҅ �"!^Vg�����g���f���8���+���{qU��<�h@x��C]�-H�`]=''��ϼ���wer��x��aT�mX�[��y�a����%r�"���˽��}.&��EP�m�;Er��#�ήȳ��>�gz�@����N��I�-Vg�OFGZv���J��*�"%:Z�-�zs�Q~�ף]��{U�Ō���8u�u��H���涄8�]�_�,D�s��Q�"Ph���ԉ�G6���4�U�_�]���u��Ntv0��"
���vB=i�j�J�d��i舝8M�т�]�$�*go];�3"�"��ݎ�h��$%����5;!��;) xh�C�'�yM�eԫ*1_���y(�K1�l���9�?�4��U����ֶ��Z�z�)�j��?Q�d)`�U�¾��K����/5/\7�L�R\;7��j���]Wx�]�K��P!��@:s�2�ț!p`�/IA$�2���@���]�Ji�'Lj�r�\�����EQ U$�v	�#��n]�� ^�\>ʥ[i��ʄc����t����9>�՜�H��}�I��t���潌�0�����	�����؈��
^8w�[��4m��##O�m��$6慳,,�&Y�۪���/�T�+A�6��D��DE�:��2M��1"����<"��E*�.��Ok�
S���c4�4u�����JU��!5?���v��_I?�Q���ZL�~������	��R���JY��%�s�ԯ�J\�������5�y�Ҕ��8���[��:��l̋1ĩ����W�f��8pŐRXv�K�^�%��C��xh��ڙ�!�N%����b��V�����qw��}a�E�d3*�|�_c���^-}�L	�+��= *(o8�%v�`�b��<��x�x���;>z�$���׌�#�(�ՠ��402I�,��.G�46~'PX�o=I����Q/P���9,���>���?,	���
�5��dYn�J�?�TKZ/�_7�e_��C�A'��~����h���&`�	�I�P@���f#Z��I���\u`�ÛU��7_#{����Ӷ[�!���
��O�=V Jܣ+ಃ�'����%���9�b��t��J��678�L��>��9�.�t
s�lM����3P5��]�<�kMM��q���5?m,Xm�u[.��d ���JImT����a��>S�j1GQ����h��n,�WV�>A�NF����[���W��ˠL��Am��cc�7�1T����y�گ���x0�!�oUN���͆0�:Ox��>�:i�</�n�%o�"\��TD���e����D�r�o�C��fGCB�-�3Hg�\��o�������)0?|�b+�"�u��M4��HSu�η�,����*X#n��׽�����-�#�E����X�8V�o�W�t�$��h��L�e٥��d;6S�J����%��m�6;Ǻg�����M�����z��l;>���C7M}����L�Ow>1�3�t�)�,�o��Z�?h��r��1��%I��E����|o4�|F��N�#~_[
pſF}!�E���ce�*��1���>4z,3�П�n{/�	��F!��s���X�3��3�f����kP&�b�d�̌`$:tk;1-���҃��C��\O���(�59���/��p����0��C{��#�ݐ����|k��2B�^��Or�"��Q�(Qm�G�8���nCD�^j��{u:=�[�O�7E�7Z:�
YܨJF�ڪHe}��+����)���o`�rg�/�o��w�fBn��jN�CL���_�᫳���	��xA�k��f9F{��1[�ߤ$���-*�C��f�D��!�$T�1w��̌B[����y�^cj]���@��R%��R�4�Y��ǜ]A|���0i`�����yړY[Ց���#-ӿb�N��l5#"&�͗�bv���ź�w��K���f$�����9K	-@nZʍjz���^>jwӷ��U��"�L~�T�P�hc�y�^��gw�E1�2誓�!ٔ�1�6:^����X��A�8R�ȆP,��D��s�J�w�P>�c���@u�&7]�h�����ּ�a�(%nu�6��эz����/�$l��YH:Qbv���Ol��i5RX����*;@i��W-P��L�n>�_�+ @:��3iH��fڸ�jJ�x���$�c����S��M�<�:��7��QU�ao��À��g\l�L�Q �*o���vȕ`~v26+�W ��1w��$�'�Pu쭷g��Ƭ�C9 B�?�uq���K�n�K[-e�k<R��xT�E�v�B?wtƢ�y���(�f'���uVu��d�ρ� e	�U�&�=�C��;J��%g�#f�
�]�pc�3�����RbnͧeZ������~��T�dsR�9	q�\����s�Q��8���+v�<�k�I:�,��\7N�/e�:�Y�K��5�#���(��N�?l��K;iv���3�0���"�+����E&�%�.�"��o�-�2���Ϩ�w_.�G�e�또e�[��_�
�'u�#]�l�:��Q&�ؚĔ�f(#���	z�C.�%t��B��'�09�c0���/��H6Q��E0�\Q�:@�R���t��d�4�Т7�X�`�P�ѱh���P^X��l��f��׬\"�F�6~L�4�kxX
�5^������X3�y�]�o>�C�I'�	B��4e)���~��GLy;� ;����Tr����Mκ����;N���8�����F`�r��+(=�a5q=��<���D4�3l�$(��U�,E\���p �?�Bt��o�%�E�2o�ɣ6M�*̂�g|d"{-�$�F���a�7�ِ{+�dA���;[���6��"(h�5I��%hHS��+(d�ήe��31_�I�$��+����`W*lE6�_q�-�b��T��5N��ɈrEA�Z ���P�;:��V����"��	Is�h�� 
��/5B�[2���B�wm�
� G{��g�)	��\���4��������zOxZ��W7���`p����o�����qw��v]f���!���߼���-&���1A�m��.���%푓�D§���執���3�����������V��ϖ�+�oy�<���!#.�*;���o���?�!�8�t;p7A�=�QB�Ф��^�����T*ڷ 56�#�� �S$��F}K�(�Y�����J�EO�����ܿ�g0g�1}̻��w���p_`�l�����f]�*M�:e;'��9u.U����4HR?�>�3y��f0�#�Lzd�jVq�l�ľ��4���/��پ�(6�	��.�����ae��Bv�"��A�^���<ٛ۱�݁y^�r��W�����+�sE�Y�8���Ծ1}՞�;-VC����;(i&�=�2�o6�����A�,�l�ܥ������}�@㝼qZ�0��Jq\��2#X�ٴ���:I��u��،	���y�b�R.٣�Q?ï��!	l S8�&����f12�iF\�/�=�ͬ��x���q})���	p�(qp�Bs>� �d�D*���f��R��]������2�5���S%!���|\G���$�I�q7/_�F(��8�۟QW�tc��¥fwNx9u��W/׻S0�3�x�
�oA0�d�W�*��*ں�hy��%}P�:&����O��$D��Fy�1OY�����]��E$�ۈ��H&kh�ut��̽�ߞ��	<"������[U����yns^\��9#�H���Ԑ����+�&�%�r�7~�J�7M�:
F���<6��;���-����B��l�6����g��{�BJf{;�D���^��S�ـ�e����h1�rE���w�S���l[�Ë~[����i\h�:6m���l^T�P��{��S]�pODK����
�o�V��S>?/o�T=Fb�Ve��f�R���.��ͩ>�c�}7{U���ݖ�����#r�R}`=�� �G\��o�o���Si�.�!��K'���ӪX<�ϥ��Q}Pu�Z\�*B���S�0���c���ߐ�(_��a\�5�� �	ƃ�e��C��xq��X)�	�m՗[eb�h�}m�c���G�$Bƪ��ęo�1.zxa��ی�p%�ѹX�O��Wu�ހW1q�`���u5�D�!��=�k��w�w�%�h6����L�$>��@�n�ŘhUX��{�8#���8�|:�.���E�L�κ��U+/��{@'j�l�1%Rq�/$"���=�'gY����ݕM��r���t��,��Ĩq��'x����ߩ�$�C���R��$��&+��(n�͜�/�1��!Ƹ�_��n�Q