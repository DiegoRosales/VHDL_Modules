XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��q���	�����I�G�J���])2�`3Gj�#�$T��7�
���I��Km(�ү8�O��4c��>��k�qK��� 	3+���̺�<L�t�4�Hy5��j�*��D��#��u���	⧻��#�9�?� ����7<H����#W�Ȇ�tv��&/' !~~j��\��S����%�"�\M\2�8�����e��K�yOC�!�(û�՜��^�y]ַ��������͊�x6}z�����c��R�W��a�J���b��ª����P���o���eP��.�¬�h����࢑$�$j�Xb��lP��9��a����hm�W���8����T�ݡ�~�������� ����p���Z@��`~䃧���to�ڕ��v`(������]�@�5R
a�l� d6^�l���H&S��)���#Q
�j����J�?,���3�n��m�LE�p18��>>J.aG���bA���+�R��uò���Ñ8CW ����h��?P�*}��L��kRa����$Hu[�]i���.�y�ؼ�����Qt�Pv�6Fh���A��9��[�@����P����$����:�L�DI%�9k(���������YC�^Ln�<�2�0��"��X�d����8�BAzO[�1��٠��7<��sݤ���X���I����4k�Lc���b>�^1P�FC��{��.#���o}m�ۘ+�7ҿ��K�@��:p�e�I�A���,T���K�?��XlxVHYEB    12e0     6b0��@�f�Rފ�\�&=;����� Ĕ�kw~g��oi���&����fbd�5-��>��,����r����ZB�v������Xm�sA�v�9}ź���H���{�bǺ�I�����@h�օ2�k�<�e���6/��F'��<�j����e�5��O�uh�@�`.����^���!"`�=�r���Yu��RG�����9��A8
�w�娿ӹ�ļ�������[l/8��"A\����:��u��f9��仫-Ғ�38$ƕH�a6!{��;g=h���U�D�f�~�$�Uu9&�C [��]�.�}�n�R������]i!OY� �H�l��!(��SQ���!�'�%2b��ll4Z	�<��G�KǕ�$�LF	���� ܊u2a
�{Q��Q��T|�h<�-��HG?_A��34�F��6��+.�t�z�5���V���@8B���?S*�gu��°6J|X@�ɞ�����L^���z{{L��9�t��Ң��̉?�v1�r�� 5�P�YL��	�Ϭ�A�Gc�[�g/�w�W��D��S�~a�����W�;����K�Xo���J���h��^ȍ��ΎĜ�{��/�=����i�� )���,�҃L��2�����ٶb'i��]����3��s��2���ěOW��:�����TK���9 �N���a�?���.3vY W��<.� �!_��[�^�<��ǯn��0�C�bN�^�qD�������b�n�J_o��[5����o����z;�v���RV�Z	��
F�f{�J�aQ�~8p�?F�ܗ��}��d��`��&O���x��V��~7ʀ��DU��/��j��&a �����2;��nE��3���3���c}ϟ�������@~�#�#�\$.|ز=c�a��+�&){p��Ş�ފ�Κ`�����4�^ٿ��=�܊���A�҈eCew��]l�o8�d��M�@EB�O��B���_���-��W�TF@'Mc�#х]�}N�������o�*�|Rn�~�V�I��
��#)���1S����s{r�G��PL�3p['I��B:�������E��k�E�e��4�����!�}�+)��(������w=cT�k���_d�E�6�X��=�-V �=G�\��X(9� %��o|�d��]����wOb[5��g$���C�P�J��D?�	'�����x�IE63���!/ݕ[��x}��r�r]���>��t������Y;�6,��Q���5�u2��b���F��l�
�� k�&�M��%��AY��L�ϻ�Ň�����V��e�����3�������k�t�}�oM�sR�8�w��Ό�ck�O�rssp$1�jP�}@痿�p=Ж�~���/��U���ŕc;��u��s�w06�W��-�a*I	�"�P��o�X�.�$?�T�gu��;u킧�LjO�#!Yd�*[�V+b�D�����y��q^�u*��O-�!��i ����1� ��z4��mԵ�g�N�������s��}��4���'N~L��f�VTУY�>dIKV�����f���G�M��)�X+f�C�e���(`�K�a</K� 3h���Y�,��V�0���W��2>j+]�)��D:I��C��*Nw��Fx�����v�\�ANAx[ʕ�O|- T5��b*��V�e���"3