XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��Sg��_���6s�E�
��ʕ�8��@X�q��w����Z���&�87��7�Br)��*�
�fX�i���J�_yB���:�JR�A�+��O.�~9�����_{f~��
��HB=C;p}uW@�l�o�����V>�l�[��j��{W�o,�=�>nk�K沎����
T�������6��٥`�Ǜn��%�!ad�;�x�A�UU%5���@E8�Z��u�����G�)��#X���rs��C�og�W�m�U�
�O��	��J�+���0&7ˑ\z��9�'Ez�'���I_-k��v��?�����D�7����<��U�P�ɓ���J���Y��]�;,��׏L����e~���4��S�f�U�뮴���'�
��]�"�o�G7�]�	"S�NΚ��?��F��{W���{~t��Y"��HUFH)�p΁gÈ�m��^vT���L�޹���,j�^~)@����{,�7�\5�?E���?��@��T����$��x�������R�߳�I�^=���%]���s��-����y�=-�Uh���~��A�w:L���P�9��ö���LΩ��Nމ��J޹ܼb̶	K�� ��]����(��%S�uݧ�FG��u�S�1ѽ*f1̟��-ĥ�bz;?Ԭ:��`�ݑ������5�+5Ԛ]�'n^KaK�#�I!|[34�Os�2����ɲK�b"�<�X�8G�u��s
��J�����3XlxVHYEB    2907     cf0io�3ެ��4A���!�����vu��]����]6�:��+�ѻ�]F��P�,օ(x�:O�]��D/�z4�%�l�/HT�w�@%v����ͷ��|j�C�3>��Q���d������=��K�� �v�t���ڷN��1�P&Dk���&W#1�O-��	$�Q��	�l���BX0Ej��W�P5�ilG''vm5��ӵ�l��C!��q���-d(g�h~l�6�KEl����yvS}ZӖY�K����t�8e��h'����;��c��qI1-e���bZ��: L͐�U,�P6��K@ʒ�=� ��ي� y+��b�YI��fQ�f~u|C�& j��W
���6]�RM���O��`G��h0�r�l��X�c�x���E\��쾤:z�#nR�־��	n��sQ�@�_&ypJt�[R�J���Ա����5�<S�ɴ�����J��S��_�n���w�O^MA��M�ch�/*U�b��{J�9}'4���{�j�ߡb�`�%#k�>s�W�����Gn�؝nXGt��No��ܾ���O[#5P�aQ�C��D�N-�^�$B�&ڢ���%eN���h.����������R}<-�����~`���;&��Fi��--C�f�X~�V�{�����9y��[��Eh�]�)������c��JD-��0&>�"Q��B� u�V\�IIr���I �vAn�--g�
���m�ּ��"҂V\|�uz�.0NRw(o�	�8:���/�	�KX�]�"`��'��l�����Zi<M�!w*K�ڏ�L����3��E���\p�0UH�&B!xU��plV���b�^�8=@��ҳs���d���l=Q(��h�2po����F�k� .��Vs �{G��?�1q��a��Xމ*��̮Ͷ{�7mC�KNw�F
��p����~� �o�����{�}E���ݖ�"&��9Ggs�����5��O녢75�2"�8I�*�W8���)޴F�jS3G4��*jTU�h�s�a����rlɽf���Y%�sK3�"�V�f8:��/4����-��[%���z�z{W]��`�I�[j�ţ��hs��������q�ӕK���N��cC��ߨ��8=yV$���(�y~�*^뫺�%_�,�j㧨��)]�ƺ܍DsR��^b�/>¸)���{d�+����?ֲrN�#�
���U�քי�Sp�dUQw��YE㛴�zr���iUqi���K�E�����	�7˦�����|!��:���ۧ� [�C�K�ݒE6Q0p�á� [�������~k^�Q�a+�ы�Py$30�'��Y7"�$ɭ��ܟ������Wg����٘c�lh�b��yQ ��uQP)�k�|����Nx�!!!!��'	Ä�s�ގ�Ǚ��F�&�I�)3���eJOű�L�	�^w���j�Oi�$�����ت�j��?I�s��b�@鍬`��E?����Ƭ��pr�0�Bd�ј~��#�q��vy�~���P�o�}�V�S7K�m�3!�K@�y��-N�71���N̰J�&8oN.~Iҥ ���(:^�>s/܂�䕶����yl��c�'4({*E��p�G��|���h�D�GA��m?~,���3����h�ؿt��v$�]�USUP'|�˩�%�#Ū1 �PB��`�I؉�\�qJ��Oa	�Y���O4O��	y����ԸD�D���}ڤ�f�1D�y뼷�(O��B8tA6��7@E�.�Pd�W���7�nb�Cf_(W;�����?�ǜ��1in:�+��C�¶�
1w���o��eQS^hѽ�:�{f��k0rӺ\�,X�(���Ș=m*�Jup��fMTI�������m)����1�ڸ�$6Mi����\�*:0�h|��2l�I�|hQ����ŏ�W��f�@�l�������Vƅ6	+o2l����j�D��^�1�1cvN�����q��H���N�|8��2x�ۡw1��0��bUrʪ.[0��E���L�ގ�vi��~ZՎˮ ��⬗PT��vZ��ð�lk�������N����-=.\�	�������0��#z8	e����Ç��٥�\���)ϲ,�	1�ǡs��Fzx�Im���4}�F]s͋�|(��p���/�r� R����ޠ5nLi���h�!;���R��-�c�4��n�4��A���%("ݡ֞.V�e?����g@�^�og[��=V����єψ΄����4���˺���2�)E���<�����o�}�ι(�b	U���c����Jk�<����k�X~����2���B�Ȳ�f�@�|)d��%+��G4z��I!��N��yJ��L"�����8�x&�AY��pԻ��7��M�*�ѨɅ�5<D@O+1X�Z�Ժքk����"�ڒ^���m� �@.S<����$Ӑ�q0�3�d�S�5����(_�Ƹ�pΣx22Z���m�:@򲪵iJǃ�p%���u���p�ӂap��)$]RhMz���"���y�v�t!�C��ό��[W�\I�`�M&7��Ƚ(i�ṷK#|���J"���T78P���Tv���8xL��nT�ox;nέ*�*���\����E�� D��>I�'�\���٧4�M�P�V�3x�L 5H;���4�������a:�;���^��A
C���2��@�i}�O�u0�[�dT��Z��%���u˵��}-O�mr�?��呅��+�CD��TX�R
|��=\�����u���QUꄶ�\h��-��׵ԛp�Rn��9�M�e&h�FV���Eֽ����R�=�"�R}3�jj�E�a��W��� �a;` ���Gz{{��PB
uN+�lԡ'��T���nAv�����Z;3G�h��ͣ�jXn��>��)�� (xۡ��kk�GJH��Gz?��o��4K������*V���{܌y�f&����epY�&���Ҍ���aT3e����<���_������yw�Kx�C�M����byɼ����jk3�n�?�����	s�Fp���=<H�D��C�-�d"F��5�%�ddsY�iiR��+P5��.�
�]�W6�m/��Ƌ����*��er��Qn�st��xta�kE�T�OZ]�y��,XW�����]fZٵ�	����N
	���XA��˩��ڤ�.x�&8�Bl�����V�:��g�1D�"ʹL�'ß�^WY8Bt�3s���>��jo�Q�