XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���Ex����MuE.�N�#���)���o��$�g6:)Z'�cc�n��x���Մz_8�4 �})��'�s��Տ'�Q���� 2Olz�j��Ks�Q(����Q�^���-���Z��U^���r9�v�����~,��l�eh90�N:�߈��^߬wFg���t{��X�aGy��n��i�d���G:����w�knu�Z)������Pvʰ��V�_�f[������Wl�}|f�D��WTL>�`�Gؠ��![`��^�$�z�t,��4�ō��P'|k�E6F�G��\�]B�Dt��-�((�h�Xr�k�~=��� ��<��#"Y�p�0���p��.�=H��[T)���M.���	&I<�d�x��g�ͭ�������e���v�` ��T����,J� o��0+E�d��]��H-G{wOۆ��*����"�2۞
�Elf�x���3��Tۿ
}���N'{�=e6z��y���q�oD�]�#�p`i�^F�ԥc=39<t��h"}Moz}�N Ƒ5��H�a~ŕ�G��%��WN�6ˁR8� 6�!��s����7=��Y񌗣;;�T�H�#�� O�ɫ��Ѩ\�3y�ů��/zz'��y\i�g�z���r�@yf5︮Œ��Iz�y�����������fi���R���T!�r=������t	sF)����1�F�
��.I��k2���������d�c2��`��i�5�BR�< �,��P��8ޘ��&[Y%��XlxVHYEB    36f5     e20�#�p��b٭��u/
�XIk������S�q9C��W�Ke��+�&�=���G��Հ��ݑ�����𒛸�S-��KCe/����W��/Ea���� �8�{�`8�1i�bԾd5�E��f5]���IT�o#�m!MWY�K��@$��ly/ƪUrdM�$���w̾j̶���8EL������	�-�ۣ�/��R�U����ŭB���ٙ���~E�=��i�1.ދ5K
������g_� 0�x�->�:��%�'�r�������|2�ϠsSiq��܂>/wa�J��������Y5+i4���6����A�(&�����"�v,=�h"�+.�@�~m�G���/�N8'dQ����\���Y(�#�MԄC�4��B��pQ��2<GV��%��I8Ze��_5Z*�#/�юTq_��l*��3OF˚���}r��l�ԂN��V��"�������#.�U��ML�;2��50�]�W�G�Kyo�)��������&�ճ�k����:��s��/._B�_�KC�K<{)�*��S�D�9���"Ҁ[ 7MA��B|� �M>�Lfѿ�k��]�5��OEi�ܙ;T���'��_�i^���� ��	fc�-\0�0����^̝h���G�ks��S����������b�HK�3�)�U��S�P�h��?����I�k ֭fM��V��$�KEG�K�0���53.�\��ܤ�²-*@o�/::���po��z�eν?��M(i
텴����Ҋ]
���l�)gy
�cmg�r�v����Ce�Uma�@t����� �f���< �8�p��#����'E���q�Lb�o�	��?",�J�
}>j�ʱ�"n�+�����s�6�{7����\�ZhW�-��X{N�,���b�� ��ˠ-/_��3��:]�zb����z��<T��ws0Aᒺ����?j��͓-��J���՚u��Wg	�+w����b�K��ц��;-l�ծ^��B���k���	Q�J �і��o���Ι��Sf?�߷.$*�?��4�^�K��3S.�P�h� ̩�����n�2H�:���f�Au# �*���>�(Ȋ�Z1fG����\�"��;��+�OFR��P� �W��,4o�y�?��Py�ȥј���yݖ�9��Qo�D�]�'#U
�g><�O�Zw �ǽ����-�0�t옴�!���7�Wd�eJ��:D�V���K�qĂd��/�}dѲ�ʼX8M��OVP����5�le����0X�����W
�X�x��k}F�8��w�m���J3}P/���������̢b�(�@
�^�/6�j����DF) 
zÈC��F	��~yS��i���=R/��7��.�|���3~{�'V�Ǿǯ�݂�M�m����἟k:�"u ^u#�yJv��Z�W��0/f��y�_M*~�m��E����Y�M��-u��L����.V�0��޸H���9~]=� �D��8I	�a#��9=0$�D�1� ����P+o򪒗�dn����q��!�_��]E����B#;j�Iv/՜�4L�÷���+ ƅճS��,�d8Yl0_K]�Y-!j1��%�;��9Y^NA�J	�z�%0�,B�@���& �V� 4���R��C��X�5?Ǘ�@�����ѳ�-�^f]K?H*cOӿ��%oMW���*.7Ym!�M�^K��~4�1c6OWq�!b"�%��{�]�p�����p5-�{#����3V^+\E�D	�y/��d5��kc�im�\\PyA��yL#A7N���G��CUX]�?wT~�_.����,7M/e�G���
hq�km~/�z]��p�V��� 6|������#�����3������rt%��Q}�g�~�_���[P�54�ͧr��� �3�=-�t�m�`$�2���X�e�f:��/6Y�W������N��#���1⟍����d��o�s���䷵�@r�9�+�ѡ;ZI�+��U��5�O����>�kǿ^@&���+�
�f��38g��	"V��|��E�~�n�z������M����u`8�./����m��SyG�(`�*U�������uw���ô}�.-���#�m��	&ȭ\Tĺʜ.՗(�g8H�w�X�N�HL>��OT�5�E}^�����T�1u�e�aAC���p=�	`�
Ţ�t`W�d
p1\8�P55�$�	p��pFti^'�t��_yk�Z'���h����3�9)Rg�����mla�+�;�O�|�j��E06"��= :u ^ܢ�J��#K��O �%�(*g<vy��%d�Y]
D-��O�(~��#��@�[d���c����i`�g�?�S?F���f�h�*B1u�7�@&��Q�����E�=b|Y����D��׹6��:�ț���N�]� ~l��)\��a��!����!(g���[Dz�i�S'�Yn�?Y(�l�|�����/8���oj���������GK���T��`z1F(��P60*[v�i���u:q�Vx�[l�(���
J�\�x�]����x	,�Um����R|՞P���~7�1&�B���o	�����P�(�>J�B�W�Й�}��l��,���,�y�Ưf�6^J�g�L![���v#/�{d��PN�)�缀V���q��8nuYE�?��Y�x�τ?mwB�1�2a��!/�%Z9Oʗ�oy��'�n�0�혻��N���ca���W��M����"�reV��&�	���{�h��C�n1c �m6�A�YY?����P��V	��[�p�����PZ�=�	�v��!w�IKZ��<)pvѫ
��-W�������NP9���J�1��S�Lz,PD�-r!�[M��N�b�]���JQE��sM���^;8;����W��QJ���Z5�Ch��N�n���}Hn%;2��]�r	���Q�Y��Ӭ����Gk��@E�Y��jh�Zn-Q��I4�D䯊��B��SH�YP��F��)���ʩ;�\(-�S2ki,|h1��{[�yQ@bS
�,���8qؙ��cb�9��Jq��T��0t������»�6n��-�3���h*R�;z0���E�+\��JX׈.��Z+��ƕfr[j��%��Esa'�OD�hm��-%���>�BM�Xx^�o̪���/L�}��>޷>J=:|X4e��9XO�ƚX9Oj��i�e^Y�1c�f�5Q�L�qK��w��"wpӢ�Y�+����R�K�̣�//�o�2��
B�Іg���H���^(I}����\�����aT�]������5I]2�C�0Ur��m5����8�Fv�����0��O�͈��������i�������g�8���
��E8��=�HM�'��><���Ä�U}�:,J'I�q��T�'S/�1�8F�N�[�%��������Ip\���C�u���;��_dg�����t'{��tHf�ϑb�+���,Eg������h1`�]AȐ��eTh^��7 �gt^�"�������o%�p��8C