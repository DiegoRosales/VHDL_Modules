XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�����-��$�ғ�i�6_��+�"\`Y�8bL����#'��\;�	{��y����t|�e-�c�$S�;��A]]`��2|+��_r���(R)FL���R}�w�c���2�7�p��l������xl�<��,�*{M�˞�*�'l�)��\��7߅���Ma����q��lvf-Ǝwn��%X����E�o ���=���F|j]�?���D���T��b�΍=�d�^��R�J�D���Y��pP�nBxD���#�;�^���_!��8�T��Xc~�u�T뫪�5
ʊU�"B�a�r^
��"čf�˾������*̳��E_tx���YΛ�]�c�~��A>�@�J�#J�����Q�F@�<����ѭ�r�0-oq{e�T_���m�L��[��ɤ$L7��eYM���1띕����97�������bJ�X���1�=a���NŨ�f��|5˴U[�L'X�>�����}APUTr��p��.pu;%�_]d�5RW`(8~�u�>��+������;������K�kD�}ǝZh�"������G�T �i'11EG�	��{�:B�Z"y::9�b��T��a֊�V �(��?���=��y�Z߾ď����ʝ�:G�ŭ��Q͙���g����T�S�ћ|��lp��u��R԰]W��M%gV�sF��_#��s�gm�1o�H�0�'߱�L�֤��aT��6��3T}��J�[��4�rB��x�|f(����o�d�c��t<�Q ��gXlxVHYEB    fa00    3120Vx�@i��L|2��·z��>Du)��Cj�A�vsyn$ۙ��K��V�R+�$`t�XT`i=��;�5�O�������u
���U[��p��rp�4G<K���lj{^�L
�M���Yfb���U�~�6�R�P`���#]�D�r���4�U��Y�b�5�?���{b���S�ЮO��Tu�7�� ��;ܨ���[�96�>�w��^";� �|$�z+��R�,U(��c�B�Ic.���&��xBJ`iÏ�5l�|�l��Z����3SA���!�
��)gG�V�m�d�F3�ֱ�Ti��ݴ~x���1?�G�H�
��B����I���>��w����xm��9C"�P9�YC|�HGbcxŴ�Ȩ_��+ r֤�<X7ה;&����&e�R�m�䈅���-��E�˴\LxF)��=~D���G��m�`�v��(l��A?7o���������Yp�65&u��8Ȅ�`���|AE���6�]�'�k�U`BSR��o4w�a��p;���k8/��<��4�Y_�X��1E+D��uc���m^�8�щA)թ�+B@g������p�/��ס8M����k��8���xT^��ffU�Ԁ�ZT� M�O���-�|�;45��΅5r]�g���(?�P����w1o'�c���z��o�o78Rha�[o���W��GP�,�3Y�!)zܑ+������zF���o�q�#vtv �8q}�&~��i�� ��&�8�j��@�Y����g��	_��R)���X�!�{�E8�s�w��T:�;�%<�	���/��Dal�VV��Yц	O,`��6��Yve(��A��7��J�2�{%'w�+uH�4�z'��6Kg��y�x�\I(��lg����K����[O�n���d�cĔ9a�Y��8ų�a��u?i;�n�R�LA��(��`g(&�p��(��t��BN�>��p�U��P��%��%_S��|X����������ɋ�Idn�@)C�	�y�Hrm�a���2n�R6�iY���2�5��e�ғ�,�ܴ.b��'tl)i��G7��2O������թBZ�R��[P�ZHĒHx�o}mՊ��a��VXW~Ŏo�Ҷ�<m-�< �2�t0&��3�#SO��#�k�kp�n�`23ͼ��(�]8LDY�~(�I�v��pA3[�V�eꃢ7�0߻1�x���~GMu��bly1E��R ˡ �/}��+q�b&��5�0�vy�ư�r�V����g����2�j��Gp�aӦǌf��P(�zĕ>q>dy*k���v�B=��s�VT}!����l�����L��![����5�ȚI��V��߅��<�|�\�~�Ov�Bv��|�Z����e���sA���+U��#���e��3-p&?,_��L q��� M�uH����Aih�BB���̤�PdUs��g�����sm�Iɏ_�$`�UR�2k7�s����RU�m4�(�A����;��.Ԏ�:T?������ܳ���r�0$0�%�����J춺��Zsg���'J���M��]��e��s��i>
6ǭߐ��0#����.���燖[J�j"�]����V����M����UÀ�K��X��f�Ż7�*�p�n�/�2����+�N���� 8Z�lӁD �z���%%����N��5 �
��T0%���Q���_4"Y�AKDn�q<�)����J;��ZiO��z���P��H���D}�~���;��\���-�u�O�V�L/�UI���k�4����e�d�8=��R�bn\|M��$�U�qK�L�"���~�VA�Q�ڸv�y����A����T�q���^G zJ�)Pb��g��iMؿ7"�jP��A�A�b��b}� 9$a��E�NAc���-���_�3�q�4�ɬ-&�'
�:��ѝ]&�.!�W���U�4�����O����\`�y����-�F)�#1��<���Oʃ�����gA�>�~JWN1���w��p~3�{VvVN�7Yy1�f�(]�Za���tXc�ѯ��J
��y%n������zӢ���ܝO�^�땅�gT�(ɟ���i���0/�Og�F�Q�h����c���"5��!EZ5�S�I_�XF�M=���#���z(�OЧ��s2VZ/���,4�w	WӱV���r�l��J��[s)6�~B�Y���4��z�_u����HG���M��1�Ј���hr9���OY`J]����8�������k�v����C{W3\�Ǎ #��E~M*���b��%(�=8��XR;NFO'(��b�s=��B7ȱ�~'���p���]wow\+���rOae�t�������D��R���k�5�7ۄ�{�;��6��dN���,�
��#3�nD�s�O�D(^�$�ݪXC}��J�[n����~6#z������Hup�zܜ����@,M蓠6��?FO%��_X���#�b�->AP=�|��4���;E*S u_�k������z��N�#u8�F�nU�z-�����]˲�=MT�*k	C��k"�t('�uNb�q�k������ʕ����!������]4�5*�a>H	���\_#mY4�~Z;g��'@;zoH�_�D�c\�I3,X�8879~�"�g&#�v��دXJa���q�]U����̥�{rrSUCG
s\����(FRt��޷�E�6A�l��}̚������Gɱp�������v����Â��� ��_c�S��>|�x*}&>��>!w�^|a��G�+�\0�꼚&���['P4	GA����iC�۴��x�{�ԛ���*I�h;��k��t��o$'x?*4yN���֬M��H�+�u�?C$�����S(��uf���p>`xߏF$��_��qC�Ł�JNr|�x�=�b�Ƨ������r
���������X�ڶ$VE��	���+�y99x#)��E���ڴ���	����c�->�˟�	�U�g��C�Ρ������
K O��/�ے��4ҫ�Q\�=%z�l?�M��;u`���q���}֣��H��'��I�3ҝD?��A����\��t�-���f�嚦�E�}�24�Vz��M�:�C���㜧C?W��a��W��X̾��xr\��۲}s�_Ȉ���8���t{���CR0Υm�y�_��d��Gda�I�E����T"-%rL�m|�%¾#�s
��=�d�-�Z�+8QǍ\F������D��~g��� 7�"��G;c^�e�J[NW�R���+gR�l�E^��3�}�����U�v�-� ?{?��20g�v�x11My(-��_;�S=��C;���|���4j�oÞ�q$K�^�n�3�,k_�[�9hΊ�8c�v�9��n�k�T��5"�������y���F�Ä�d�v5��B��h��t4j�1\�_�M�UM�n�������L�>1�]��Ǡ��`(��)��;#��B~�O��4o+h�l-Wa��}�ѓ��R��Ω8�MZ"� <�ʝ�A:��x���c$��v�ND��t��S��	������#G��X��6X�������s�G5���(P���)�?l���@x�-/�*�2����P��.��-Z*���)j���d��p/����m���Mh_�����Z9�	�I��&o�1��'����>W�$g��f��g ��+��֚ ��A�K�'����?y�|W~��2�����%��ƴ�D:�˔�Lb|H�L�9�HB�O�`F�[W�}�VcgUon`ls�-񊵇zѺ���0*�Z v+������L����=fm�C`�`�+'X��c�+���5K���p�������X�q�R���I�^�]Y��T<+S��s��>�m�}{��揉�}�0�@���p�M�D�����2��12Ad�_Q�t�G�i=�9����:�u?<�q���*-���.�V&���z"�s':�h60<=��Q��F�����Bp�8��M�Q8m�tE�e1����
���dz��T�u���r����W/q(�'��/p
��8�}���o�UE)�e���?�ߥ'�A��R��� �IB���K�/^��}FU��hk��<M��2NF��VϥX�n7�@@c7v�Y�,@̝q.
�KÖ���+<�LӁF�����,P>�nI�!e������ �����L��Q���	���c��W�@r���zIM��k
�1f3瀋���)�!�چ�� M�����E"��k̍�P��������g�(��g����Ao 9��5;�m`f����nT<uYA1�w6[	��{��֎_<��ŭ��h�L��\q<�׬�H�-l�٢��R��_�7�*uW�S���Wˣ5��s���$ᘥ�;���c_=\+RyΉQO���j����WwM���+m(��R�eD��L�zu
:D�K��� �[_N�Q��p��/q��@`4���F�$Hz�?:���G����c���G�ص�O�S��s08��w-�U�%�/퐔����'����"��$oM�U�jd��2e������\!qF���9�XUkp�u��D����:�˜Ը�Ѥ7	����Ꮖ<&�l�K�m{�/��31�WY&�hqڱa��,��I������>o����N��`�W��!��"(�AC@È\:Tc�:������{-!�LgE�?e)����튎��d}2�]�͚��F��p�9���~բ]9-��&�'�Q� XÔ!�t�*��X��K�m��&�w7����\+�%���P��1�H/᳙�Ξ@�n�@i��7�p,�$�5+�{h��[i��q�ǀ�����c�?���q������ 3�Rwu
תB���m�������Dc^�p�	ě���Bu�U���}�0��0[ C%�#Jȯʂ��N�l���D�
���6���upra2p�)�;�Qi:?5�B/!���dQ�fI\�@v���A0��G��i���)�0�L5�K��	�V[���|!H��-��BhV��y4�S��'pM>����|��^W��~OT�G�$!����C?���ޛ����3�A�VO=KE{���Ɯ��j,�KL`�
�/����E;�����CD�>����5?u�܂���>�xg0� ��Y}Cn���^��A��֬x�x�ӌ?0vՀI�xH�e�W�U?z��!�^e:ÿ'T7Ԛ��wA�f�i�	!�*���@���g����j5��b��أ0iz`W��1�� n�]5x�Qq���҅�..7k�����R~���K{s���_\��E(�B�7	�A+=G���,�DY�5x,*�.���w3M*����5�s���O])z��/t|��kh�qV9���J����5�aRp�nɝ����(݉�D3$G�+�T&�hJ8޺X^)��c����P����6 ����s_qz�th�A�'��/�̠(_G��"3?,���u]N�5yt暀޿��[A�E�Ԅ+m�=�A��Se�����>�����-h�]��G̉?g�N�v ܠ�E:��#���B�OTWU\��ͷ�qL^5S<�
f�JC��B�Z��	,E���\Б���� �+��b���7Ⱥ�S���@'����f�3�J�c>��L.�ʤ�����@g�&D��v�а6Wy�L�%�C�?��� u�);'~T6�[�w6�PeR����:$����^�X½
UJ���`ȻN4�4&?��'���m�V,1����珈L���Z��u%��JH)�6�_t 6�_Y�wÁ��0�A	�ظ6����e=j�.�+N��/I��`~1���D�%��N�t!Iz�נK=��� ?�(��-���|����T��i�dژ��MQ@bO���w���Q������U����'F��IJ�a%{��0e���5�g0�QT�>�F_��?��¦7T��y"��>��1,�Rl��d%q��5D�7�Y���O����E����|$����Gb�|הte	|����̼�DEz7ؤ;L�O��'m����L� �'J�|�3��>>����5N�f�-�o GC_$����1�E�+���8I#��_5� �"V*��d'.�@[| >A�t,��Wf/��pU����ʸ+�O�bsvg˝P�'EFQ��^�rZ���jF(c/Y��'��7�L�̿�3�&���~���T�J��
�K����e�:rd���U�>���TPp4�0�S5Y�����*JW���X��,����/�穁K�����ك��/�����?��e��7�USr�&�uﳄ�uEn�戛0�������%��M������_	@�G���0��<lh��G�wXst9L��_[wF��%��y=��{a��.S�2Ĳi;I�d�%���/B��%:�Ķ�O(��s�L�~?U͆*T\�o[������m��}[^�U3���l-d�����{vHR+��Nqp��f�i��N������G�s�X����<�l�[4���ִ��˄�J��^S�|q����S�Q'���Ԁ�2ym��G�9�kK��a3@W�ޙ�Z"վ�&��:+ZxQ�Ddeg�R[�Δ�Lh��i�Y@�zC�&��裔���RP��mxc�� +(�kV��J�K�uj^�8��� �߰D�����*&�1 �%2Xu���;𔡏:�#���(���� �o&�_�Fѐ1�O�]`y���׃��� X8�<��-���U�Ħ}�fq:��!��E`L�.h������n4�{m9S{G�k�+=�Y{�{d=�h��1�ǣM����Sz�����Gն��ٳmAk�W
��۸϶|^�z��-b/��-l���.$�&�pk��nmm�ۈ�����a�M��'�i�"
�>�J�h�	��O��6ƲBk�o�WgE�s���������79��2#$�6? ���0�}��Ҫ�tP�\P`I�,�ڈT�0���"rX��oC._$)Xak]-T�\z�����2�����U8���9�k�H9�4�(^� &�˲FWa7�!�e#яr$
�	|�"i��L����R��:B{j�נ�+OU�{�#�k݅���?t� -ߌ?j\�d푧ԅ�+�a��K��Q��aXά�D���"d�y6���
� ,aϾJ$)�8���9^�s�`sc�4���ZL�@�h�3m�!�:�t�v�[L>`q�����I
@�sۉO���њľ<,��k>-�}AS��R���2�����(�e��G����Bٽ>�|�+E�1���i���UX[7�խ��� ��2̺D�l���P<�U�\;ر�m�ɰ�w�HISȨ"u��|{�(��C�7(��!D�x; ��_�S&!��"�D�V�"�f,�Ҥ�JL�E�#�܂i�:5�_U�����\$r�R0t��G����>T�Gr���k���Üof��l�Bv4��=.	�yL��܌�������>�tI!N�!r�u8@h��j��^9٧+BU@��8�,�m|�5�/����q���ՄL��� KB�Ͷ�ŭ��؞A�����qW ���� p��{�8�����=� �����/5�f}쐒V�_Km��P!��Ce<l����~`��O�3�c�{g���&�v����`�Ǽ���~�偰�5>b�BF��}���������U���.�1�ޗ�G�w�
їE�����v�,pφ�)?������ջ����TnB�ޙ�ӟ��X����S�����>�zq��
��HG�+�ϲ#��ʒ�I?c�?c���9D��M��"pA�/M�7̼�i.��i�,��g���$�{Lf�Z���L�?���P=�gb���`�T�r�ޮ��^�L�_m}�F�uc)���$��vU��n�B��ϵ�au�l�:���Z�M;�(�
��"K.ѫ��Mv��pq�N����z��I�V��j`	��q4zk�##ܡ|��� qK��)�s�$0���v��4�_&�o�U���j<tjHl�>�!��2��s�7��aIŴa�L�������<B�+ʮ؜�4�A�o� ���ZE1!�(*�8�ڂZ��Cl�ߨNZi��t�c*���.m�SEV��)F)g1�jm�m.!r��ؔB�0ƫl�쁺�L�0k���m�t��2�b��W;C�1ROQ�m�(u-���ұ�R��h���z6}v0��JZo
���o�u�!촞��>�x��f���,��}�G������c��|f>�E�آ;�Q�[O(����`�ˊT��,��(�%�Ѡ���L@B;(�Gϲ(�*���0jXa�@jr��K���q�M=Z�9�������}c�kHӶ<pʢ.�~LZ�u�y�3V{Y <r2�`�.���kv��R,���9�k<%�a�bk�n%��<�~71Z�]���n<fM�_fq3��`��"a��>Δ�A���>��`��II�A��Y��U��$y���o�y-`�%�d�8�b��j��� "�< �{,޴�j���/|�� 0m��\մR#�����L?/J�!�\ZXt�]���`�<5�	�j���ܟi�b � ��� �	148���|����'� ��B^J�s��d��&����@�<>�s��bʪxm�q{b*���ڏKM�^qJq^��?�J����J�J,�h'�e�n�d�[�b�!�j��Z��	���1�f��lY���K�I����4�_�b�h��,CҖqJe`Տy�b_֤UC���ĖQ(����"�U>J��%�����B<I��]����9P�]�İ�߉'J_����3�n$|�54�$}	Ѻ�"{��P:
j��&�F�֕-��y^]���Q��|��+���(�#L�&L~B����2�
�)P ��Z�
*�7 �a#�6�s�s�g�9�(�F�}�Ja�CT�P�%�k&���x�4b�7��1��hzD���n���@sQ-�۬ �&�sU�Ȝ��kB�U�[K̶�`d��IYT�lMj�8\V��f��_�4b2R� ���O%�|&S�N�p��{)�O/���0��?bc� 0gE��|���i�qh��HU-�оs!5��˶V��E�-�0�B��bXv�_�AG������׹'��.�E*���=�����c�,�������5o�#b�U�w)��y�=�T��3o�ڥh����li!{�����	D=�-$ւ����&t-�Ĕgg�HT|E�LV�[c���xY��7�5{����ٝY�� �J��Ž�3NT<j�=�G	ܤ�+��{fSZί��?�8ݲ��>�Q��)�~J���ͤJB���f��� ��w��]�������*�
<�kS��^��g���/R�W]A�����>W>�yt6��
��g�C�����RK����'Gh�cki)m�(�|�p�����g1Y��:qA�CD�������c�)V��/������?�\> [����2� �������R.O�Şݽx�s02��V�g;*ʯO㫬�x �~�O��Xa�DҊ�kR�fO��Ww��~
5��{t�Z��FPY�B,�%�V����?+�7=����z�_6k����o0�i�|$$N����z|i�9=�<��v#���ebE]��5����Q��
Hʭ�����T���[��yt.��8�\	B!�N�dY2�Q)�>��˄���l��Mq�>���(��lJ����D��Y�χ�︫�f���UDP��o|�,�5��.�%G��PaT���`�a �K��-�UĤ�#�������[x"��M1'�+U2݃އe�:JX�-�ez;tW-bEtPA^�1�L��"QEgN-�okҕ# -֬&���mj�B&:Z�2��W��E�G�ز�bA9�̫zt��&L\��F�>�J�I�4�c�ht1�$ ���/0Y���8ᣮpa�7 b7nSwX���գ��ٖc-X-��v"A7�����-�����X���vf����Y���q��|����2V/Tt�?�z7����Ȓ�7s��N�o  �S[D��#�pJ���&fy�	�=�>�2�JRPFN.�03(���嗚��	!	M'�F�-�RhNŀ�i\Y!�a��x"7�8ʄ'��́����+�ѫ�9�u]��H�g\�;��������n����@�-�f��ҴZ*xb���k��Y'@�I�,@ C�������0��g��4Y�cT�ʹ��Q`>��U}za�~�D���ZӒV@g��kFm�M���u*������޼��- ��Zj�:޴A�܋�u?���j-^f~�����[Q�B ;^Sl���
D���$T���W��|3ځ���0�����}�ߢ�5�����'2 �������[4Y�,>���ܳ4�0C_H��@	�c�"���n��c�AC�JTࣹI���;���G�X����N�!���5b�!�<���H�f�v>�����h+��Yf� k*Z�`:&@!�Ɵ��������	���e�~6���(S�~� �Ř�q}���O�wH�c8eiLڌ��4ʥ���eXDȷm����`�v/7�'���K�ham�37��U��r�R
2�}ZZ�Vvl~P������`�盛}zp��򣹘C�7��f��5Uk���ZM�j����J�%ɝ�3�rE�j�ge���X�xɎ��o�m�����V��Y>d. ^o���'q|�J�b��NOx ;�JIJ�r��q�t!�������+���`U�խ���jZ�y�M�iG���I�K�l�H?@�Ʊ���toj�o��xV^�RF�o�8�|�2?*,��H3o��[a���{�7AU�s�?��h+��#��� I�?�+���SP .vλtW�&l��
l�$�{�&:3����p� �u�1r�+D��,�E������k�2��j��k�fZ������z�^��JpX!���%��-�|.�}���O,*h(x�u�ȁ�\I�K���%ۮBa�3QS~��+�aQ�߰�s�G;�����Y���_�X���\TP��l��|{�Zn��Ī�a4�3f�:\�v��".�G	��j�h���&�D��� ���e�1�\�Ja')x����\��$���҄�x�B�5,�ҭooI65���i�i2��B��U� 
����W)�h�5��-添LES����Uw�y��Qm�n��H��j���Y�Zz��JN����vK:N� �8����}7�K��"���D^����˱V�ӱ��P`�I���¢������lU{���h67�j��D�-zF��!,���f\��'�v�	�ci���s�]�\�qCD�ܧR5d`���t�4���$^f�S�BA�N60��E�����u��sM��
�hɠǕemi�ޟ}���ě%�r��q�Q�n��EE���ŵ3���
OQ���1^<�Yl��*W��!�@#9�]J�b�� ��]Zb͢}
�x�r��d$���$�����6����t�Jʷ��s�qTR!�$�S��G���L�FnA���:P��N l!b²����i�G��4�^7l�;N����(\�'Of��eM>�V؄@�I���}	�Gh�2�ar�s(z�1wO�R�����'����!�:��ǻJJ0rv(��0D��κ��^����J�yl�F{@.S�b-�4zB�&��X��zA���3�dKyX���gQuj�fR.'KK8S�;~�y��*4�TE���p�sh��!��9��#�Ʃb�n��3�U=���da!R� �Ubb�:c�F�lpA�D�˝����qU~��4�������c���g���,�O�Ӷ�w(�i%r0	t<Y��Ty�����1F2<"��;<����a�nmu�jꢃ���(�7��g�g�_�Sa
�@�}�|���H�����j��l"Ef�����0(o.��`�ksx	Q�D�#�j�������;y�pyIo����l<{�������I�Ga��:�\�y`
O֮�Q[�a�G�Q�\ڷY�b���#�e/3$�	��i�F��\B����zN�HS9�z�l��}���S��y��F�������D8:�-XLmU`qFJ��u����s&��Nm(z��˥��9W��V��x�xo>�@�ZG��C�϶�p'p}�j�п��=��BFՅ�H<��r�ꎼ�����Ed|j���~ ~I�
� �M��P�{vq�C����j,�k�0l1ELg8�|`
����K3�YGc;�Ή�W��3�e��� ;����Eބ���f��kC`t������9�ܿ_������+>X)9�3կ�%Q��mAq�zV®z��w�Z7���0�6S꒬Y�}����^���XlxVHYEB    2311     980���nk'�-ؗ;I/��m��F�P��4�){>���إ>!H�pP�f��6���ow�AMĊ��բ�3j� �L���6<��2"NR���o7��쐡�\
�^��ȣ΁U[�v�X�)/6c�~�������ԩ�r|1��{Gg����3(D`�}�uh�z����(�R�=i�@N�><O6CyQ_MeW�ϴa~�ŁBI��QB�>��y%>��	8U�{{ d�2�a���,� ��q*1�sx�;8�v�~�'��vCʒ,VQl[�|������4�r	�ӍM���"��V��خ*��b'M��vT`�'�y�)H��'�Zj���aw����=w�L��s~�����'T���u��g(ݓ������e�X<��8�H+��۶U���9�#=�@���*�c�hn��b*v}b�m}���7��~��Cc�	�q׾pGK���9�h�)��;��Mx��c%�|������� ԩ�(�<|����?�'��H{���F��1��2��Hxi��W6�dVRLO$���\�n�߯F��D�c��﫬�#������e)z$���D�`� ق���B��@gG�Ǫ��#(ŉ�/]��bп��k@wʮEލ��<��W
W!2��}Dc�y��uM�lN�e�Y�fU��~d�䈶.ȿ���ً�0����m|�ڲ�H �;+������~ݯ��੯-H0Ot��6�3���!">uS����f<Èa7*�tg},E���P�9DT�/�\t�?<�'�1Vȅ��ޥS��2�St�"�+齶��i9h@����f����Hv�d�{���=
�>T)@̈H�&��bc(��i�|P�)���뎧H��V�|Hͱ�F�S1�
f��}!�X_�"����eH��bG�~�����?�վlً�κ�1�PmΉ0�p�����Kx���0Q����k�p�P����Rj�}�G�$h�\�ڈ�ڗ�.��eG�J�C���%����ﮪ aWq���ԣ�=O"嶷�7���V�p�^�p4�D�dͯ�r��A �ޤ��oI�L�( ��b�~\g�(�A|#F����kI�ze,�/�ҘW�@/3�l�I�:1��"va+ñ�Wֵ�X����;	9�8�hE�*�b"+_�=��HyDmןS��O��Ud^c`(Ȉ�z�j�k������7�ݓ�+{�z�v�"�*ӑkX&���yW���cY?���2����>.;���\憿:���/�'�:�_Ü��p���e��ܫ��P��w�����V��X�����,�r�}ߤ�O$Ջ��<�s1;L������-4��x;����w�E�i��5ƥ�6�[>jo
pT�u�xHGKt&Ӝ0u�%��ؤb���(��H��x�ҿ$`ZY�EH�&d�^5~�zˡ�Vݙu�>!{(�ʬL���������P�iKӝ��^��4< �.	7�O"�'�}���>�K��%,��M�?������f��o>�8~�L�ɣF���u?Ꟈ_Z��Vύ`�lR���;�9�1�W>tqσO_{i�&�I	����D�?��K&��Ji�7��������@�&\ʷ��$ er��R��<��-�<�w���{�?�J���'z	"g��1p���6尯�����d
@���������K�~h�9Sgy���K���h!1�qJ+�Zܦאs1��k�tZW�N��p���͛�
�� �y�j�"og �O�Eu�GDH�3T�w��yԾH���R��v+Bl茯UO7u����g5
z��RV�i1z4���\j&��ǜ�M�H���F-I�bTRW�90�л��3�/����ܜ�3��`�E�4���^��h"s8��{�Z�}I`�q�Eup��z�}��S9ō<׻��mJm��Y���L�q�E�G>�7+�S����Y�c�~�[E���zO6��@%͎b9��z��Y��I��c�����W5-��$˒Sd�����궫?����$�*�J�<jqS�t�X���� �����Js8����t{i��3$�
'Ӷ�=5����y=�^<���ڿ?*�th��Hѵ��c�vMN A`�2�W^tâ���,�ȓ�y��/b��{N��>��c�J��k�LnW��%!B�k�G�&���Z5;�K�u�^������dZ��� �2�z[n�zD�LR �e�o�B�ƺh�L��&�*��1i!�vo���<m�e����8k�qc��4��&��S�O�ht�%I����F�>WZY���M�n�D�9�+�#����D�
~e��`�"GI}&s�S����.k:�J���h�d,����΄RH����:pn�p��\����H�=o�6iC�ټ_��I�4�X�&�:�A�d�{h�����