XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��O0"|s���B	�Vi:u���y!ٻ�WArNg�E�ތV./�4�@�Q��!��Ҍ�-�nz|�uh+�~E��MIg#)��4S�w`|ږ�"�6�S2B��j;� b� �����Vc����F��9r�V,���4�)җ���%%^��B�8�Z	9��d`+_�d#��2jR)8�	�<P�0��]�C9���:����P;AMsU$hL�[Bm�J ��V�:�sX�z!Ymu̬F�J�P�E%
~1<���<�b(��<[ ��ZD|cJ6Ě�$L�49%��֜���\]��g����\!�
�����  �ό\�/��W�̉�}\Yq&��Klj��cQ%K�F��ģ8��0twW jp-��2��y���-x��xG����f���x��8�Vm�(�[c�e���f:��e�٣��@N��`�XhŜ����͟3<���V�4��?�OH��3�����\܄�Dϣ�?{�����!�g~���0�k�BW��e����.d|:�>u�. #�4dqV���3|G��1����x���ǵ����t,�h���]�
h%*�z85�7�l�Μ$TFu�,E�,���Q����]��m1��M�� *��cF J�)_�Ւ�%�͉�T�ڝ&\h+�ȟ�}�3��w���Q�z" � �ȟB�@�����{�A��M�]Û�$i��� ]��d[XO����e�d�8oS���*���o�j�ӑ//��!4<Z!�n�j�D[!����XL��XlxVHYEB    2163     980kT�����%m�h0s�J����(MO��d��������N���!4�׀%�.�fݐW��m_ZR���O�%�jaIiD@p-3�X;�q0R&�P>GD)'g__��qk6�	(Nu_KU��W���9Ww�{P�:��B�\��Q2ll#���̧+�'B%?�>����3D���ٴ2t ��j*��D)̈$�YGI+ȧ4�w�m���Q�A�\9��2�V�z}�&-a:�jn�r|�?fAdi��>{�������mF�U�XDyIPb���M��+�]"�+�'�^�4(�-���|��!�YZ��8U%���/����\2G�s*UQL�e+U&զ�DT�$Fԗ�f�a��Q��Oc��w.���K�܎n�A~.z��Z�<��'w,o��������̤ �}�uC��ֹ������7��S���|�ttؤ �\;1J�Cts��������^�W�$'"uĳEXp��6��kG@8;��P� z�vP�9��P)t�9����fs�ү/w��L���C{*`�}`�-]�-�\J7�I�X�:�F�'=�k���f w�񦙛���:�Ж�ϊ��.�>��L���䦷��C?��N*��E?
�S秺`��K�w|�J�KC�/!�[@� � �\���t�\Wԇ� ��}�1ۓa.	�F����Z�8J�hй���S�m��Kaϙ8�O_x�bЕ������B��U��RP�+Þ�a�K,�W�L��7q�� �����_�mܚ
��w����0�!_?��6�Y�g�G��������WrοYF�������%����_f�-�sUbf&��G�=u���4i��t�_֨�]�����%�7>��<F�6&6�`53�
��p^nQyp],e�J,-�Z�@�wqP:��5˷��((?��v*V<[`#�(�b�[�%�:*��|ڳyt'�3�[K�z	d|jqe*>� �W�2Kv!�	r<��$&`�*��"�(�V����:�e����b��*�z3��q��ߍ�o��[�د;���j/D��8�7ƻ��y�'Ž<!���3�%-�G�釽h��Pw$�5w�ɺ?��9�]��m��w= L�+?s6�e$Ǡ�Brbv����M���As}���бY������2���Z���*�ힺ���_���D�+�/0���%����sa5N���
��k�"d�=P��C�����v��ۿ(&�4x��J7�|9h�a
�P�pk��S�h�N։�f��l�&!�v?Ŵ��^Db��4�)�d�.X;�b0�@/�2�&�9��圕�R��-�;�b�� ���W7��;Q7L��)r��C�'n�F%����B�Ι�W���.y��r|4��S�9���n����T�]c����R��J�	�����C�~���$ץ޶���ͨ^�h��r���X�ͭ'T�ٶ�:�j�p�!�T_�L��N�.��5t�%��)��s��V.:-M����<Kj�Dm�o��>74�y���6ft�i�Ҟmm�V��Q�i~����M}&����o�[rk9�����JFY3Ί��Rϸ����J~3"�+K�B�hdS�h��|p���'Fqn֞�$pA�i�=�elR�/�uϘ�ZM����Ȱ���$[�{7��k�E�@�.*�R׵�p恹��Il�4[����������$v�d�y��X.��@���L��<��O�;��'B��bHI"�iU�����U�lF���'����`�.��Ճ
�z�#����'l2&���i��Ә����k��$�~(��1�,Q/a��3m�H���j�}��#�)RR�ep��9�l��$����]���I 2F��P3�ζFC�'������� X���gj(U��.�8R�yI��O?����+ K��/�i��Xs�i�s��&o�P&VqgehJ�]hY������o�qǤ��==g*}Y�)M�ie�vi�����@��2�۶~�)sC�����0x��!ޔ��`b�ēu*�!_������z�#��ڦ�$�H٢,<o�w5���L9E\���	)sXa��b�x���� ��y͟�H�R�X�R�����M%X~�4M��T%���ȟq��r9^����%�������C��L�*��0��Y��P�V��@��6��ꔏ��;]����ϓ�K���{�D]��J�.M Ō�{�i�O�b�b��ZY�U��d��'d�����N�Dy��#�d��'x-�����Y�i����yr�4P��fg��)tVӗ�5�IBs��W.4�t�E���Tg~Ș��a�jc	�IC�]��L}�m,�r*�H,ۍ�1�]�� fV��D��kfPPГ���
� '�7 ���Ã׺���U�oҧ�|�"������H?�