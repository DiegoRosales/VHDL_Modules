XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��3�_N�γ4�Xmm�r�g,�8�|��9�xŰ�)�b������®��l/K�y������/��	@���B��\�>W�FƟ���L*"��[;���^���x[l�qw�x ��F�3��X|���&tP�^��jF#}>m�6�;�.�@�@+=�K�\��LO�	F��a�_tZ��  :�lGՅ}�����Pf��1%���f[���[3nPH5�qMs�=��?@��#��i��8ܬ�o�Bg��Y�΅�F���EbYv�Fz>;1&J����Δ�mfsL{�+w�3�̷hR���I�Ѿ�%�:ũ���5,#��g�	@r���V+S�g���dՉ�Q���9��8V �����!����X�����Ȁ����(�Z�W�"t���$�A:����pl�X =�,y�)�8d��,B�m�4º�����U6Q��c8��n*�p�k�/%��1`[�V���)�Obm�+.��h����|���b`t��K�H�A�ɲ�$��܌Rg���Ddf�8���V�oɐdK�!�n�Q/��������ɋ��O��gL�娂��_-hj���y�l�����/�
Zh6����/�����D9���I�T%�
-4��`�� b����@��K��L�o���sG�X�xᾇb2�"E��u�L1�H/a=	��GK4��}�A��v5}ќ�L^��ځ
�?�_ ��v){�zF�U�@U`4�`�+�����[^�T��Ckj�}��-_�8��w��0ܬXlxVHYEB    2447     ad0{T'�~5[����^y�7_���v����>��vY��k�v��8�zj�Vc�榋��D�b:켉pT�7�]�,�Ѣ�������1^���W>i�k�V�}W<��_���-QSi'2�m��Ǽ�@d=�9[���.�,���Ҝ�O����+��<���:҅�%p�����.[���eP�[��n���ʪ��+����VE���چ�m�7j��L�:��^�}2�	��gi���S���#�M��1t��풄;��tO��Z B�!V��f�P:�%K
�L��O5�o����u����=,��!o���+�K"S�t�D:-��S�W�0������N�1����Z����ü���}�����$`�r����� �o$K��7U����
�<�?��������R��A�W�uE�Q�\����O����fL��(�:�薮���Q�ꌳ� �u�벶?F4��ɝn�3?�h}��ʂe]���Nj��`J�`��]Dk�����	~YL���l���b)!<��+��ΰ]+lMT�'D=���j[�H��bN�Dm�ӗÊM�t�kkB����� ?T���⚋cc�XA%���v�(��ET5��K\�n%z692�n.z٩��>y��+��b��*A�jS�I�G�^�_8�H���?R�)�gj�ܧE$�^�3D�@Z� ���Ey
� �\����
L�M��SS{�_;@|ݲy����52y�|�i��@av���WBmn��:�S���WV�� ܫ�z�=Ry$��tr��W��q�d��bgRk��G�cj�_y}t�Ѝ���C8��㑤y者���z�ކ-��̾����h�|�G�u�l�S���"dG���G4B�	튢��7��^���̾yo�9>�O����P��� ��7�=?�;�.���VQ/����~�6���=�>p�Fu��o��T)�8��"�_6o��O
�O������F;�?f�c=��M�5��9O[-ޟV�{�	�U���ʻ��\��2 yʦ^2DCI=�|B��H�D��R�c��-�?�[�s���"�]�Z2�@�3��|,m��(/⸿�(�F�����I�~O�ѡA-F+���n�11֖��mZ��`]呼��<J9ӟ,#<��ؕ`� ���AVK����?0���K����S1C�'����X3�!i�G�7�o�:[�}����i��שS4��lٱ�1����k��.GAܳw�1��ﮎ	�'9�#�l�47C=���?���֑�)YC�j��;R8e郤	���v]ȴ��7�����)�"���k������)=�/�����o9��Գ�C1��a�E�4`9O]��K|o��U��s\Hf�5XBݎ�݅<�D�@\r�=��n��������ԉK�:s����e����x��_�AhTL���:�P�&e�W!)\i�/A�m8��)�
6I���cs�]��Kd�]���a��I�"��'T�� `S�*-��}+�&�7W��������H�,���ֈs8�(j�j�1P���L]dX�:�o���黅��u͹�������f✈߫)� X�v�ܞ�u����OǇ�Ժ�>��6"Ν��:*R,�d-it�³V&�5��{b�ȕ$0K�0;`��#"�����T��u����\/L�#�yꈫ+��w�|b������~����p�l��a[y&Y�ټ��&0��苈rQ]�PkG�3���Y�eT���@&�=׀���s�:��|Z^x�'�,�1`+�%;V����AmҜ1��d4J�'�5���ɜc�8s��d�)�~
�wc�/�>@Xx'�������3��I���r��+�j�{DE%׋�#��|�PJ�+=S�^�m:�B�U�U(mv^d3fP��m	���U}3�@��<U���5��(�|4�V.P�L��	�5���6����y>]c�.Ҧ�)gw��^��,�T	PX+3�UL߼D<�[9U���%:	�\eC����|70��$:�%� V�q���'/��s/�'0�j-jd.g(�z�������"��:�/̴����T��Oh0O$�����uHZ3@�A��ǜǆ��V\�r�O�n<Ď�C]T����@Wj&e�`6r���	_T2Y��L��܃,a�N�!n�{���e��c6xm86�BU'O�Zc��1>��\�d���j�)���A���o�*�P�!�#]66bN����k�vQp���韘	��)���^��'\������>�?jS)�G��A���M��;^,#.-O���J�8X Q���k"�Ҷ^�c��>k4�ʴv6u����ZA?K��]ׯLӆ�r�e�sC�9��8�\ ׶"���������$f��~��n����2&?�I�)�ώ��X!��is�Me��<W���B-ү����Sl�|πi@�\ �F?�O�t��:�ow�ǄrqsW��&���|X�$+L3�_���k�2-�\ϑ�)�{�Q���f�a9š��CD��ŏ��Q�/�4"t��5�;m�����t�&{��m��ǹ+��;$ݫ>�L+��lޡ��f��éM����?���9rFCɘS��n(��~�8���c�rL[�P�Uk�$ ґh,�1�X��<����ׯo�t\�^_��w�-W��b~�8$����<�e�A�Qc8�:���������#M��1.�whE�흆2i�σ�j~�