XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��B��3�?l�s���2�)�\��(�ٖ�B�m1�H�ŖK� M힮Չ��cW����؏yR20����.��m7�^��^K���ޥ�D�����zjio��6�Ɛ�J�U��#��9�����@"K�nJ�Mh!�|c��!�	pFe��}���!-�y,v8��un���WwO���l� P�6�����K���^5)�T8���iE�K�Z����7e�Hǻmn�2�c�����Vҩͣs�o=:�5�l�HN,6;�h,�g!]�1�RړU�e�V$�΀YVg�����G�S��SV���b:�e�aW>ᡮ�V��pԊF�,��̬'�t S�A�����]e��-54��Bʖ��w���6�	:��k��C�Cp��3Ita��"���bI:O��er	,�u��u�Y��w<�����A Т��B�{���<6��a-+��%�.T�2p��]���~�띮t�X���ނ0+t�L~��9��ӑ�xҕ͎��2���y��t!�U�ha t�(>��9�]_�4���!����Y-��Z��)�	7-ׂ����
t�G��j��_-�g#���)�����{,�)�MhU�ҷ�G�\�c_�&6e��l��?S p�-w��K��	7�"b��U�A����f"���Qa�{��P�V�ٗ����P�T�o��W�GKTx當uA����j�*,������+�B����IA�K��L�(b��,C�P�fF�n=���s���B��"XlxVHYEB    36c2     ec0?��Fj�p$	q�&�0-��]#[�lW�������<{,F���<6�ힴ��$�f!Z��Ɛ2�+������VS��AW��Q�7�ݾ4�<��cav�OF.�����/]���i�%mp�D�#G(�k��q�si���l�,���{�T���{	��evun\�Щ;���ؖa��B/�͒��_w�L����NX�xïa�Cbӷ��;�"~�����>�S��,�i\����ӗ� ~p0Wscy�Ө�9a,Q�i�!먀+4	/��}����Yjt'p�:�}v��{�殀�������e����i(M�Oo������m`kDA��O��5C��G�yQQ'L#ma���fH�x��G�[�p󑻺�]�*�5ݗ�� |����X�V����{�:���e&�1���u;w�ֲG|���>�:Ŕ-yҮz����q����Ű�pGmp� �}Q:�K�Щ+�H�%���o�an��DG��*�[�m{���ի���g�' �G+O��'��Ĳ-=������G�rR�l��JU�`����e� ��b��6xo�v,Lfa�㏍şU��x0���%�f*o�<|0�P�Ǳ�<���U|����7��q���]�LY�pT3{�#���:��Q]�o8��9����ޖo?��b(��O�y�j�a���^�&g���),� s�|'eS�S��l�܈[A��d�穝2��]����pz�G������B�EX��O��섀��!O0�RM:-�7�FAmzh��G|�%^ aU�j	�_�d�'�$��(fOAh9���K��_|~��>�C�{�陸l�.R�	h�c�x&���1��8�s�5�E�<[�K"���$�bem����e/$Z����ީ$�^HT�4�����$ ޿N:��w�Z{�7$=����鼓�q�V�+!��qw�!:GIݿ��C�nJ��f$�Ul i_K9 *0sጵ84���)+]ž���YNtY�����H����_z��.���͐?��\�%��j��)�Y���A�&���OE]���]HB�J�oZ��#̱@�ė�y˘��R|F@�7�o��ib��`�85��]6���o�؄�Ѽ�9W��P�mT��R�2嫿���s��ċ�c*���D-G�����.䗿� ��,V����,�L�m��TĀ���J��&:��(�����	Θj�cx{���ԟ�-#	��~ۆǗG�W ������������FY`�!����S��`��A2�̳�#fE���J��o�X�l��L�.L�	Cd/�^~�1ꈂ�"kSO0_5��OQ�o�c
����`�,�I��xq6%Py�q�[CO��׼x[zv�u �YE��Cl잢�5!�`E�m�0뒳d �Z����p�/�"pE����yfgVp#1�m�{p&^m�d ���5�������g��r&��T��^~��O�ߧ�NɄ�E�����X&ʸ�Q���{��UG����w=wq5Q�pr��?�AEMjȓ��#���| {-�=�� ��q�.ȭ
�`_ޕ6�ꂍز�G�2�ݒ��.���ol��O��s��=q��/H�@Qp��@8��{���"��7_ë��)]U���%-�%B�"�|���,��ۓ(
�L�I}^gL88E��ӿ����ۧNPkE@T@�;(8'.z�t�	��OH�X���o+�~U����B��M�<L�[�n'܏��6�
p�w1��8tA����E�!\β�����xd FR`j��Z{'�b��N�ە���ٿ��+{�y���ј4�cA	�29נ�~�9,�5����I��ǻ�|ڷ*�b�븯�]x�ON��(�y_\X�������ׁB5}ř�2��(a��r�2{��`�,�,��U>m���'/�ҏ��7��ʉ�����3�ЌQ��Sͤ�@̞^4H�|"y�?r� TO{����&�,YeL�{,H����ʌq�&��j�����5�����5��F	`|Co٩ݽ�`�ҦL(����N��4nNulj�2��#/�㠶�Ŵr�&C䈎�«��)��I3��.R̀x-�Û����A�C(�������0QkC����+i[�������5vrt�[wĐ�m�h��>��S���YZB8�;e���S�f�F�JT ���;4��g8�$��:��ڦ��OR���mr����Y�2U����ok;��i����X��g�-����N��!JRw�D�	�ɟ�b�ss'��g�<����$@Ͷ�g���`��=�QF�͐#��J$&
&�17�
�~�3��|�'�oX��h@���e�0n�\L��`e�$��%B����8O��I	���Tz�n��7��}�����Ծa������9�������Cu���-��&c�{`N���
h�+\�B��/�j���=Y�`=/U.6�H��`����_��UG����V]��=>�Jr,�&K���)�b�_de����$�uJ�WQ8�z|l��{���S�M��T�3����6$��8��і�$�>V�y��I�T��~t|�. W�j[����Uߚ���8�Vs��E��֥�Y�ȴ:X<�'z9���B�t�#8v �~4�ص:mOJg҄���c�H��?�g�����7 �I�Y�=3ql��H#\c��T�B��K��a���.��ƐraZ�p���д�-��+����*�9u�q�2E�o��}=D�0�*eFw�b������^�(�Q��������Cj���.��~-S(���Ͱ�3+�M�0�V�����	:���̘�UZ'��c����Z���Ct�:��7��J�JW_�")�*�5�A@��v����b.+
�bPU��Sh����=)�$'ҍ��{��>��Ͻ^���P6Y�y�y�͓#�7�Ք&�'��7��!�-�U�?z��ق�b|
? ]>S�2�N��+���	p����vK�@H?�T�]�^�e1"R�&b�,T��VC��Sa?��E�3B�y����[�E�3���&�=:i����d���jd#�H,���a�/?u���r����J� ����w'w;"se�G����њWc��
�캛��'�{�ғ�M�=БK����"���M{���sʎ��e�gZ6�ӝgm��}�V�>!�x�z[&�i����#.)R$g���Mͻc�[��|�/�σ�2 ��3��MUu���z��{�"�V��"�{	&��u2<_�N@��[u�Q���y�J�Xj�\��D�L�N�� �	��3U��f ��.A���W��}s�@����H�u(���>K�,ҞZ-|�G���)E�{`r�C��"G�ns��KP�?T'�)m�G.�M�v/譚�0���x�a?#���X��.C?N�����4e�y�-CX�ˑ���F�W���pDΫ ԓL��<P���I��u�Z�\w�P�R����OM�����A��}M�+��4YSez{�iy~Xi;��z==�WH�:>�##��-'@�f�:�A�w�i�P��e@J,w��j�S2�ʐvC�۾�BH��ؠ�Ԣb^��6s�ÓBl䠁棇(�Ǣ��o=4�8�F9?���a���%J\{�e_�u2O�o��N:soJ�c8aZ�-Y�xjT���+E_�^�~�JІ�=�;Vy�8ǚO�M�jV%�U�j넱$C��Eǽ�f����(�S�;LՄ���&��\�L��"��Iv��̝��%%�r