XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���/礥�"E�}r����m��� ��	̏�0����ĐȘjC�<M92�dN>˲�	iB�T���!�cL�/ݖ��i<�㤜�9q1�o�&���W[.�`o���]�
��ʼ��{j��u�Ԣo&�˳�ɛe	��S��aˮ=�����D����Kj�׌/Ĕ�	��q3��w	JgB�B>͛��33������'�z�۲u�Ubՙ;dKQ2���������S6�9�� *5�d�`���H`��P�!Y����� �[v!�
�܍c�Q�P���Y��)�☚��I���쇯f�\�4���L�R���ʳ�[�CLw�,�Ҵ&�ƀ��N��Jj�aX�FP�E� ���:��ﺏ�M�.mWs���&�Yeq}�J
�ȟط����B�A]j+��[�h8��L'L��SJ�����6��?��In�Yy~R)�@�ɶ��O4�{A<I��ֲ>)7�63��y&��.3��Ȟ�F{Z4����2�NF}/ݷ�	#-e.`���(z.�^�1�����ԫ�0�hSwu�_SR�KV��A�Es�82����Y�^�Å2m���C���Ғ���El�=��bK���%�[t'��y�0io�m㼤�B��X��Оg��q8�����Y��AoqR19I�%��}	$�t:�t�uIJ�~����_�(�d�KS�뉑V����U|��{V��N��#��@ 0�a� q��J�<z*���'��-��XlxVHYEB    22a1     9b0F���f@��7 ]�����LT�6����4_����i����5�X@����{ɶ����2�׻i�QM�1u�<�����aH�1�:���H�>*�S��ԏ�.~1[�b|t���u��t�
 ��	��ؚ+������M
��	�'��ߖy*�`��Q��-�ҧOtK7%D�g�����9�D�3c	Gm�8����mhV��]6 ���$[�q��l7%��O��;�1p�>8A���z.�IA����/H {����eE�+�Eag��`��jQ��$@�mK��<�ѻ7���.�ȬG�.��ק�a\7C2�f�M����������2Ɋ�rRr>��E
#��p%�S)\��>>}י����P���JN=n��`��;?F���G����m��=^���Ods��l�q����	�we�;���7�%#3^TXzO!4g��46t�}=�=7�3:ٱ�%�kjO)�&	Vm}L	�c�w�nؖ�θn��M&�{e�d%}��oƓ��!����%L�<��U�n�F_T��
5>�|i����p��l��w�P.�[�����=�Y���g{��-5M�?łP�;���t�uA��u+����B+A�$L4�*^�YE��O,���$��}d�����j���9dB�y�i7D������:�(ڣ}G"�OOтW�C$��ܿ�<yu�k�@�8�"EW&��8m_>zׅ~r7B�%�+԰1�[6G�9h>�|T��w��1��U�i�-z�����fn�~@&!	Zw>w�O_�l���7D�z��B`&]x�Y����a`�@���Ǽh��e�L��}|�0���Mٟ���(��Xu8`���|�C�	TH�F����˳t��9D=r3:L�w�˧�SО�m���C��:���^sz^g���na&�S�xο���-��Mؑ��v��d��K��SY����k0)JY�ڱ&�l��[�i�w ���卍���_��oh߈bZ򰂊���2+ˑy��#�S���<�ZeV�
�v^���W9�^ֈ�0��ё*��z
@�6ֵ_�L�,��f�b��1�-y�i�]P���V�	�{,�U�x>�RU�4��3�e��_D��iWd����D�B�T��>GA%����<WQS�m׮Hy��r�}�X�qP���?�s<.e���|����y����Ӯ�r��_���(��.r7$�f�
��o*��9�<�T5�u(����)�c8�>��T����@��w�镧�:Bg�ʢ�h�f�q�O���!����B���z�br�Ҭ(y�-�I�;���Q��^�T(IBȕ�j�y|o���B.�Y�i��X����j��m2o��H8Ň����J�BW��`#�����'P$��oӱ�!RƄ��M�������Q�qѐk��x������x���Qt�݉�B���@*҅�,�jVd�S	��f#=�L�-y��Rܮq��É�M����ɘIBe�y{�������\e��!1�A�#��ղ3�a�P2�X���E��tf�z�q<1Me��9cXqr-{d։�u��L�����ƐՊ��g����*�����EEJt��,ߖ�,jx?X��|�4)X
t�>h���/o8�?K?}��q��,g��6	Q�#�X��3DS���i�g��ꌬI��Jџ���ux��H"����If�3�QǇ���OE�!T-*���2���b��
+f�l�N:��x���j`��E�o�z=ܯ�V���R��J~�ē$�ׄ�sƷ0��y[v�B�G�<��;�]����������1�gr��jN�Jf�x�X}!�KD�=+=w{
;���r��z���tw$����j�U���Wm_S�e ��`�K�����\]��CGd*�Z�h��Jj��Z�]�)�8��/����"%���$�r[�>��͗l`e�*7Y��2�`׸uV�D��!Q�J{���]髲���T%\����>�m��$�G�	�\���fs���@�#�z琚v"M�������1��]�p��DO�T��nB̭G�ؿ�'��g3�Ci�w��ʮZKEL7�j�F67W�:��"ro"�:�xƿ�w ��r�:���X�~{\g�@���/=��.�7b�i(*`�J���g�[_ϑ�D���"��B?TZ�a�.�M��q����9� C/��q�(�k���r1�7�PS��$���`i��A��^���:
���UP�1H݅�(�HD �{����t�[�X|�W��	Z�����U���0��r8U�Kқ���)�,�i��-jI���Hr,�8�� Sw���.{��,�r��^Uy���4׿��m�	��,ި4׭�x��C1��C���K���z��A	<$�P��� �E��h�!6G7��]�8=��im