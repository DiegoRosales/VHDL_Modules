XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��� $<ۭ5�&� ���eϋ0�ܺ8!������T�a��BP������g'��eY�vX��#�TrQ�Ea��r&2Q0>���pʤӷ+4��� #��
��i�<vV���T)z��,��[�O�Yb&��ǲ6F;4��Gц�^�O+b1����;&7h�:�����.u�����0�	ې;��)���p`�ZQ��֮k��ǲK�:):�!οC�/S:;�BI�;q-����B������h��h,ĸg���i4�-�!o���h��5:���;Ȫ���oV�XlT[*j�T?�o�� ��#�@�bU�)���+�aTG̚��}ݨAbI#���	�+��kݏB�p'tO7M��z$���N�@S�m͸��X�_���G<yzj�S1/�'`��;%6��)�z|��e������rG�i�br�T))��όc�.�5�e��WF`��y��m�x��0Ӣ�!���0FI�����l9�
r�)�>_�Yg%u��x��9dR�/�N2���Zs�\��%�������|"�2���m���D�y�: _�ՁA��#�ų ��	cyOqX��"̾�P�$�����m�W����q`�fʄ�i��C;��<œ*��\bA��Kl�S����R��}z�G<��~7ڕG�u�m��r\<wQ�N&R�~�)gM��ZZ1aQ�2_�YJy������?g`{�sT�֨�$�P���>7��+��8��IpǷ+%fƤ�q5���N�|�ND�:e�y��g7�\�^�X����7�XlxVHYEB     97f     290�b[|��E ����� ��_��bݖ������͎����ew�{a���fwBd��+�T���H'Э�iYUA�� ���݃0�P�t���A��#R�8�9Ƚw�t 9T�����{b�?zqk���i���͏��?�uz@�[@.�#� ���}ɒ�X�i������OY��MDf�x!vw���a���R�x��b�e7�y�@��ɐ,���������ܫê_��n#�?-4t��#�U��͆jy#A!���ڎ+��t��r0���� C��F��g�"�����F��w���J�e�݉~�Xz�]��x����'��Eۏ�V?Ad���-�k�1�t��>�*Ő�b�f����R��ՙ�6��{�?`c�lFh����ܿn������ !��d��*[>=��E���ns�;�x��MIX K�,�0�/B�&�7���Uk�<�++����Ҕa�a���S�����l�7+y2N�\MW�q�&�FZvM <�ozo:�Y�XWLf���%{���S�/X���~u�=��;@�N9	�L�F<G��d� ����ts7�(�%"ұ� ��>?�dU9[�.ǘ��!��)����՛J(zW�R|~���!��.��˥/VI��w�drw�M6l��="��o�#�4��6