XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���CCR>'�0IGm��ޘ�]f.��'�f�v_c� ��ϸW����;K��P��{s���7[�?1��|�fr���7�	�"z(��t�bU�8�7��w�kį؟�1i� B�������6�9�it㑉���#�UW��R}u�]�_���Ik�$0�bs�r��Q��Vu�����l�� '-	�S#��l.���Q#�K:�ѷ	H` 2T��9�sҨ&lF�i2��6�(����H�ߕ�d��!&��qx�?�_�ƚ' _1}��;���?�tA��K�����|�a�9�!�b�B��&f�/��6*X.��(h��G;�?�n ����	��j�o�x�qlYt�%�j����a�n�� ��aj�q�&YB;�޳��a+�2̪D\륱���d�o*�MF0m�v��� f�f,�L�F��0fB�i��ء�m��.DK��dH��&N�!(�?[Q�*���^��>v-��߁p>}%��A{��l+�׎-m�tH���!��Ь��%;����Q�N5i&�_��T\HYW���e�.y�j 8ɨܝ��N�(�/k؁���Մ��"�hR�٦ܬ1�Ѵ���������O���Y���Δ�N|�I(
��/OH}|��� (9p����-y�Ј*���&z�F�cd-�4X:h§|_/b��)�����WUc�D;��a*��^�:�٪}�үr ��2lL�>�߻
Ւ`��Dnew�Fj^)q-�)c��!�hZ�|��(X��>��ô�M�XlxVHYEB    175c     780�^��!�r�N��D��>F�{��R=Y��8�� ��'�Y���dd�ݱ���Y�V��	�E��w�Sd/�B��l���!��eoͻ<`ִb�29PJeZ�vD�7���@n���Iٹstwj�����aX���g���Ja���SWWq@ǁ�eʒ��\֫�}�� �E�C�ZWGM�Vx��A��T�
c1HY�2E�F���������h*z�Z�7m��j�6z���N�:��x7����X&aR�fz���2q����/Q"Ȕ�%�^ٕI�>&XK�Ê#Jo"l0LHϐџ��e��v���y��wT��O��r|�E�^a.:~*u�g9F@�[��Y�s���\%��=�Ep�XU�7V��"�jЖ��vr	��߯�EZ���X�W"o�Ri5��~8����/@		S�G^�X�垄=�7�,��Q��-�Y�����#��&�yQz5GS+��LqB������ƽ⓺�<���4�7����+ư n��Hq&0Y�+��̸��ʳ���?�Z�]vGޑ�����M�j��t���qV<P7|�!�����k�|
V2L�
nk9��?�u7��� ���A�^rY�K�V��p�m��9�O%2�_���}�����n1�w�J2�:�
ǆ�G,s�i�}�����;�F���%�����L	dx�5�����qmn(��T��
�C�K�C^�2}Ыy>�3ju�PghP�"��-��М���&�hٱ���h�K"D����ZkO�1�i��W��N�A����E�z�oD����h�M�]��ep��?o�o��;AL�Xh����ug�Q�/���N�C��B\j������*�T&��b��%�`����d�<����J�9(�}7�΂Rv�w���*P�Q!C��fdZ�|^������?*�`����'ں4�e��a���F':�a�Y�PD��!S�0z�K�g�tGK�?�$|���P��*��]K9 4��%)�H�r���HW�|�_Wg�R�ܣ�j�nR��ۋw�Q�,t��2� �ZHr�x�^5#��_s� �5����Hj�fSN�f��*+����fy�f�I���J��V5��L��Àټ���ќ���m�`$��&s�-�(�2h.��cyEb^�S�;��s� D�0#���VBnE�00j��	��5x)]�~Դ�<aZ�ظ;����`�fU�{g����>�p� 5�/Ę��%/ Y���	8��uݯ�E��%v���(��f������d#*�M!j�ϫ_9�]Naj�`��QZ7 w�sҡ֬~ �4vc�EU���M�cz� �5"A� ���X2�Y��hb3�t�(fMԧx4��Ñ�_&g6\lS�O-kj��F�S�H#�U~�M�t��[ T�8FnN�P/}5:�_k�.��9}8��b��s���-�t�&ئ[��?4bkd(H���b���JU������7u�KaVN��@Q�юYH_�=����	>�Mf�s�'dXjA��v
`���7!��G=��'���L-.����F��vc&j��yY�#� ��!4>ӽ��F/R���d]�����k����2��z��N',�,+����ts�n��c�_��u~FG�A2�6S�t	������>���-�hgg�@�v	�2n�T��=^F��`.<��0��>�G�ؾT6Ь:[|N�i��������v�
�	4���,�������4l}۹ůL{�1l��; x�X���+��h�%�exX�eHF�o�A�����o�$�*�y&O9�wf����Χ��a"NU.��SK�T�M�^�{�i��dz�s}Y ���դh�|3(��lg�_�J�.#�9��i���I��.k9���$��ޢD��h��0��h8g��D�͕|1�7FPCl