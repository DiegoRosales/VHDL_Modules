XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��&�տ�r����|����O�wP.��;n�-���ݐu{&��W��7�DƂ�Tv����E�?�)��b����p��p��b��4��B�̜��cV36�y�c� ��l����_��U�u��W�Z����TI, "��g���w�����b�=.��X��Jt�b�.̌�/w2��]x�3Щ�kd�SZ��⢛��=����;8WssL��~����&�ﺒ�a8�����}�kC=UB�}끥L���	���J$Q����y�� oB`��F�q�3��:���t��\�r$j��<�p���C���+����.���ٍ��dkӈcA[L�I�Qa��󠭙�d����Xx����!�ݵ�{������f�'����}���ˀ��a��5�_�ټ
$�`�6p�.��txJf��z�z�zm+��]~?(����E��o;�j��L���\���&���0��	t�`$�����#�v��	�`�u��d��vGd)5*��eɶ]Z������1+���+�j�f�A����Қ��wϡ��;w�&��c�6����;Ƴx�~���7�ƿY�P$g�f!N7��Р��9�$�(vQ��Ϻ���$�c=��	 0fo��B_�$^����g��X{<�Yf��x7��ɯ9�%�7����g��_�8��cwڣ]�{���t�SE�����:<��-��h+U��1X
^�_�������iA~j�@�?~:;�P�HR��P�_=�����(���XlxVHYEB    17ee     730���HgaB�G+K�@G�Ң�ͭ-0�&��đC=\�:,dc�����������W�~�3\#{:�E�[v���룷�Sh�l��ʡp{�.p��9���|�ˉN�3z)��r��`�?��,[H\��c����pF�߃Q�>��l�+��yC4��r��2$)]Ӵ|!4SoJ���\&�W��P@U(�^�=u;!����H����QBJ,h�N%C�9����k3Lf�?c0U���bK+.Nl���6��'��F���3R�dF�Ҧ��G�HI��_�Í�jV�r�f�ǜݎ���@�<������\�e��.�c�Jb�n!(phyo`�Kj�V�w������d�͔BW4x��66C�ҭ�RT����&��VN|�l�
x�v*��fÓg��J[�(@Y65�l�^����Y��^��q���F��ݡS�#�dl_3�"�-�;e�NA8\�d�u���4�Ta}��1��Q�)ɑ��S <o�}��־yr ��K�R�����D#���o�}�J9�f�2}T�ks���ot��2�	��f #`:��t���f��6q\6�b*��(��Y̱;q#���n��MLh�M���Q0?�7>���,C���J�*���lG"*x1&�z����D��?ӡ}>b����p=!���=:�	*5��"�xzڗ�o����*Q	� �M3���T0\!�)�~�7��~@R�e�Iz�A�@�c����PtO��)�H2�d})��V-�R,7r�0��Ұc��"��,.����pE�W��14��gϣCv9l��!.Irڵ5�ӊ�}C��6B<�����7�ƕ2���˸�X?��ι�o���r��}vFᰏ<r����U�*CĮ]TNkZ�mtH�.'+�i�����4�~`X���P���Y�~4�V����m�qZ�L����}(��e����/�j4����{2�V��Ԡ0j�\��]�y��Y�˷L���Lx�yƒ���Vu����U�G���O�0�O�v���`���Gg��d�`'@�(��K�"�l �59��N��ǘ)�o.��{f"�qy!p�q�~�\������)�6!JN��P�$�֫=��dN���H��V�^�E�i(
Tm+/W��6/�Z�����O��Xh�ͯ���_��r�*��=x5���U{M�so��k-��s���߾�q��2�!�|��'E�a�L��J�X˴�&������L�]�19c1^4��0Fl���/��{/zg9�����ID����qy9�և�yiN�UŐA�(�:��@�%;//�א�����9T���{b	h���d�O�rEIvR�.��Zn_4���ߵ���mo2p%W�Q�`�\3<;R|��3ꉀ���
��� ����w���*"�=�r�>촑-q�"���>�ʹ�(�����G쏒qƛ��TH�V�1����Ɨ>��>
$j 
D�� L[~�6-N�i�`(h�l�m�$�E&n�=F�����$�h(�!����%]M��ײ���e|w0�(㫘�� %
���̣�rik+㠾���6�ꊮ��c����A�I��F0���o�~��^��&^������Q�e@:{+�Dr�׾`f�?�Z��
�`���١�Nw��LB��O��_�?^Nn܉�I���Ժ��#s澪�S�s�����4�K�����DY�����p��h�w��Iq���Ásp�Η��������:����&���eܬ� �؊�J����CB^ON�뵠BM+�,��v=��32s��f��˩�oc!��/E]M3��q�:chiA�MbH