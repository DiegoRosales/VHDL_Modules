XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���	�3KKz5`�Fa�'�'Qw&�i�<XcņX^߸y�Rt�X	�E�`p�U�����Kɚ�)U��tEU���Қh��U&�^꾿��M���%B�Nȯ�_E�����VT�����f\�bm��uk���8B�~���?�&�3�<��u	<G"���D��\��
����A��s�:�9��#r�ʶ&��456o��7����h8��Ѩ��b��=�����2%>Id[�w����12��(�E�����8�(f�n��?�;�sZ%%:��6��H�`$�UEp�R�|v��g�$�� �:���c�ٛ�N���߹�H��kͮ�)�lD�{��<4��eJ^Y�9���$H�T�� ��D���\�����@L��cE�2pz�,b
�A>8�Q���1�*�)K`_�^��:�q���B��I����)s�D���!�ʴ����`��=FKE�����6��}u�_�H������F<ѷ�*�ޠ�^��ꑛ/sƒ �lu�N������]5�m�:���g�^Kv@��w�֡7	��x��f�n�1�k�e-e�tl0\�L%��Q�1�&�!7��@v�/3�:Tf6y%u�֋�����$���!��z|U�}����S]aA�T4���aV_��T�w$Ʌh����8�3�w$�6v!��R����s��u��D[�N�c�ocS��2��n~�?�	�o�M���|���
5�0�<idI�����<��[�6k���}0%�Y�t XlxVHYEB    fa00    25f0��Ja�\ř�>>�I���@����ʚb�M�~���?����!\f��h!�*�"���{5C�`�0����d�'ُ��d�;|�$�,dlƹ�sX~(��q��C񨪢��N���fS�柬K��L}�Z�yzUb6e����C}1����A!ad�w�Q T�ˣY��,��ցDT}��r@�&{��4���vu���BKU��lGH�pwU2��c���G����ٖb�2����7{��"D�s���Z�[������0�:�WZi�_{Z� ��c �Ei9IG׊��`hX���rD��
��ǐ��eT��ӂ���/ҕ�=��$v�IuP�&�7.:�V�"��t��9�Kx�3�2	�k�5�x�����(hP,衠��=7ь�)��zA�0 k���7�+p]���ղ07���o�����+`�-���y��0u��~��)��4�{�������B�n�a��Q{�J�Ô����L�ڊU��]��K7�6��ׄ�0�y��l7GUX�|J)@�T�t@2uܶ�}y��'�4��Y�0�GLA��fr���.�����u(�	'@����	�A	sI�w\pެٻ����)��ߦO���%�촾�X�r��?�ed�{�q7c FO����WF�����<=��?A���3$Rg��v��K�na���C%�B��yq��a_9������I��9V��"��l��2Gd��uٮ��q%4��7.Q���J~iC�a�r6�R\�^���%Q~P#/<B��U~�Q��x�e�>I�Al֪:ݥ5��2f�N��>Q�~�_\��;��p$1ww�4�a�����
�*S�!o��X��RWT��u�Jt���<&,��ao�.��������ST�eI�t[�lR�v�O�4עymi�=�v���N��2�:�Օ0��dqL�WFN�Z���c�P������:׋�ު�-E ��̅����L���,X��m|�v�٨�pjGȥ���2��8�ƥvS�ԡ�\�Y�Jh_����'i{����{;[�T���Q�@���Om�$��5XUZ���Jd�W�ɦ�o�bLcH��k�`�@͔J�f�s�Ӌ0~� �-y��X�䝷V3$@����(�n�{/!`tszX��j�Os�l�\"�]�|!���1��zX�� _����FoT"�Aė�����&Ds#��`(��:�9�:�-����|	[�}z�}�a�L�O�Ue�_ё��ak�O2��ic�z�"7��d� )������c�Y&�A���:^G~p��	!Gejc�ز�b� ��U<�ں��l���ֺ$��rm��$/]U�mL��(�3Ì��	A�����=2�\<��U95QX�I����E��滥��,�[P p���<����h2'
��A#a[A6��X;�ծ�9�H�:���nX���օ��gCp{��0ޜ���y&̼A�4�+����OSVr�r�7��M��0:��H�Q��25>����	�[�XRJ@�q������L�k�L�@��:^C��:������e�yɡ,�]�&~�dQ�,"��E����ә�}8Ot纄��*_�	�"�4ge�ATd>SW���9��+������a\�'����8^��g�^���p�;�t���EWM"2/�]�B4���ڋ������Ư+R�J���T�.��LTz�f,�� ����fTV���֨�����f�x7��)���P�/4S�d�������(\�s�����3������ᎏ���m��8�%�U�'�T��e�f�U��7���|�7@�[f$'�A5�C�)�08�|��k"� ���Oi��e��W�?s�7�$7�8+>����uS�O��Ɔxʭ�\a���*a�o>;�a~ϝ�0+�l����{��P��M_�n�q�_�\'��?}���Ywy�$�Wvbs,RE\#(�{��Ķj?�K�$��~���a��r0w;Lq�ӧ%�?@(��w�TaT�{�!��e��n��>X1�3�Gk1�����\�ʎ��-Uwj��@��#�0����^�o&��qj���f.��b�Jj0�.���<�4d���p���8��S9�,��h\)����堍h���t�]<���@��A�L�����q����擹t\�|�%�UJ�q�T��&��]r�$�YɊc�x�n�`C:� *�"�!�m}hG�,�Jt��������:p4�J5�D�$��
��臗�Gp�B�������x#�����B�p��2���^+%u�z:!��a#�Q�.
���E�ˎ��; *wai��}YH�`�an���q�⯏���0�R.�rR���uº�Z��N��Ǘ�רj���_8�bfQ�6��ck��S�Q+8����4����/E]�'��i)`�t���7����I�Qm���a�%
��֮6}����[yJ\���nL�����C]c콐!�/���2]�8�z�����
|�9��B�ݺp�����Ҡ����I.���(Q�2T�����^�	�@�*@Y��mO�&�t�d�և��@�>ϥ��ظ5��}\��\���Vm/^.JY��
��=���f����F�u�>x��l�q���d�©ދj9�r��.�{����]l�e�A"���6|h�m+����; ȣe�C�I�!�8�P����D�k��%�Z1��a~��D�oS�Ν��`����$��׎�@mHd��u{h�*U���=���tQ�W e<�_�>q+5��\�3��<�1�w����ㅁd+c�?�5i4I#�
�������$j�2%�AH���~��@@(|� .,��7H��t�ST�"!���z��W�yu=�gh �,Y�B���ؚd�8�����F�W I�%X��]PҬx�����hR k��f��W�Ո�nOe��p�j�i��	w��X�3���켪�c�,
t���!��E�#��×ܯ�b_\?�Q�3<@Z�O��O���z�'(+#T%:¯�X������z������eͭS�7���:,�~�X��	|���(1]��'�N�T}� ��括fB[�6��QCW?qu��;�~Ό}B�
[dQE Jp�q���jv!�nWO����|�dx���$z�cw���y�ȗ$Y���x0�!Ͳ���ܸ�J��	�[�O{�߮3��fi.,���V����-p_�����c<Ȯq��aV��ߙ�ǰ&4V���w-V �m��#߾| si!�Ll�w�Ik�1����c�RZ�[�?�O�[����^ď_�AY	��x����n���ti�C"��:����������@�����ZD5NC�ک�aϺ�����~�3xm(���Ƈ�{nZ��ak�2ldl��R[�{1��A)��lpy7;�aٍ��\x�pnP�
�T�<s�@�Ԍm[�ʒ5�fs��m��U��id�J�1�>����w�<�B�ϐgj�g�/�=�iƳr�n�J>�:��L��,��(E���òs��8t|��*b��j�ҷ�C�Rag  {m��{�;�������a:�} ����}�8�r[�����z|42e����OO�+��G��eX��e`����Rɏ-�M�Ϣ�ImxE��"ZѼN����i�X�z�~ѡ�]5f �n޷b����`L�����.�Fb��s���F�)�����[��u�%j���d�i?U�.@,!6�[�l�,��}k\�7��	�������u�������/�I>&����=���׬�0@�\�;��Sz�˒�_��Gy�=�� �ͪ����ǰ~C��[����/;�Q��J����g1�@g��4(s���(���#����(�L&Մɕ奚r�{�h�m>$U	#$N4+����q�َ��c�}�v/���x�'����,j�5!1��ġ��'li//��D��GU�����ݚ�M=�� ��lܰY��e�f����Rc����2���
p-��A��tP�s�|�_��l����"r;fz΁|q��������
�$߭3�'��D��'4���PMz����� ���2&�r�i��h���ݎ���Uz��_��8��mO̽u���2�_e�ͫ�Mcy{Z�j'�!R-<�"L>Z�Rz�]��%7��Щ�E�ԡ2w� 5�%_���>GY�
��B�]�G�Z>z��W���N�g�d�D1�S�_*|wJ�t$t�:�gq*y'�=>�6�ġ˄��B�}TL�C�2h��w�D��>�3U�F��Brg}��� ��@��� �Pks����7�ޜ)Z<���ɖ�=ލ��,�nng9����A�ڙ��Ϊo�D_t�-��>�DIUoh�n̬��A�6�+��)���Mk7yGtߺƴSʯWX��9�XNx���e�|7��̖��f4 �`Of����izy�To�s��S��$�#R�����$@��A�"Ş��SQ Ljy�B��l>^�J�4�o4���-Y�R���pvZ�`p��8��4y�R�d�?=��ا�������Rk��׮p��z���bd-�^�.��z�P!�q��#I�s�����hI�T����(�U����BК�fb`�����蝼?3�Z�f)�R��@��<I�ގ���� p+&�,Ro��e��M���l�o�C��JJ{��D����u	�*�}b�O)�!,;�H����c���`������ �=����9B���O�X���k��LG�O3�(��5�)����s�	zӇꤡh�B����B�����;#t�6���-����i��Ϣz�C�2�>����қ�X�H�e�Sm��N�mܙy�Y��>BT��(��Y)
�l⎤F��#��/&M퉩�q��뺧�}�g��.����EE�W[8��v���L݌�0�z���J|_k-ܶ�]��|]���F �	�qp���j�r�> z�:���A�ˢ���(�����̃��yE&�nCL^ј\��D�$'f�R�L;�������1	]���fO�q�ѵ���J�|y����уD��Mp:��88���N�U�1�.��`����i�@�b�]9���/�}��J�H��*\{�"��,���ɥ�}��o�Q�����O�4�N� �4z�{{V8�绵�/.R�G;Ѣ�*�"�"��ť@�SX�ju����1��&�\� B�*�ӓ�%����r���A;��T&�3�8�QjS�v�Ps|�#�m���Mן�`�-86���G2����؎C��r�0���n�!6�9�O-�ߌ���EC-���;��RLp�cB�jFf1��޽����;	�\Hh0RU�aQy.�i�6����H�wD�ﭵTڔ���w�52:�.[Cczo����A�rx�a�J���(rB�1�_�8�9G7ܻ�h}_�����}�u %&Y�4"���� ���HH��J~�:@
(���~D���/��.:���x�0~���O�5Mͫ/���R$(�>0)� ��4\4.�� P��GrhT���j;���Yd0��64�u����p��ѻe~��.}]h����(��8_����E�³��^�}��	�;gP�y핍�O��2�P��W-���@�(���*z2�e�����Z��J�]$��j�=R4��͉��.�E�jL�E:\K��g`��~Lk���]���ckY���F��:�����h*�"��׿�j�g{˥�&|q'��CV�10Ŗ����3H��X��MNZ(��W��Ǎ������`�:,;L/��&�x��?�����e�1��&��r���5���'
b���ğ�*�\fg))��X^�/o��F��(\T���CS�t&7�$�Af�!�,Y�,u�.�`��H��-�ʰ���S'rn��7��M��G360�ۜ�fɔw3�C�������Od�FX���v�<2b�N�M"ڧ;&r$���A1A಺��-�k�e���ȩm�-���t�g��;��������6�v$���#���g;5�Ւ�n`�򑠞��>DI�R���j���&��V�#�2Z��S�o�I)�X�R��X� �c��U��A���:G���d�O�
��P�ݑd�#-%�U����9�I�u�S�W��Ȩh�
q��>�500��r��@��19oUuBï踡3����ϴu��U}��m<4zaK��d�[�H�@7���n����-�ct]���Hz�A���a�^�{�C��DDqh�i�֗p��9��1*m)Z��	 ��s%ln�k��o'�_K����T��G�H�'��:��D���K��
'ұ�<���o�U��<BpN���9�:L�l�X�S/�R�tX����^MqRNǟTxV��~�0YS��������i��G��@��My6��}׋��gz)�n�K��VA� u���E�����U�	��N�g�^:��}F=b1�aNA-.�R#�d|���,��,��s��{
�q�ӌ����QI�Vl%�nz��ىf�C���G>��Z����R�)P��^��d�:%�y�$�	�JB��'�`:>�� ��q�������Ge�+#����%�(,�ޓ��:s|9�均l�� �kA�T ģ]���7�$Orָ8e�ZKX��Y/�G<t�s�7��3�eC+F!{�}Hndz� ������O��75��2Ø���p�JT\�ݞp02ԧ2�
ܵ����ٙʍ�صNL�گ�8ӱru����{y��Qy�<��ӚD�����R�HË]�; �M	���\uR���	��&�D6;��)��Z]qzQ}3���k-�v�)pFP,T?���S�Q�v�EN�g����E����r ��\���7�)G[��q��]�,�4��Ff��\A��ֆ5=���X���ތ��Ng��7"�"F����A6���uL��"�2�_i��K�o
����6�j�����W5�E�D���DͼB�E����ћ\ x����H�Fv�����Vvb1b�d0ya��z��ڊ��7�` ��������K!�:�[bJ��!%_fw�?��<'�|tZ�:��Lenʔ�����X��y��(�I��A�Ļ6���x fEVO���f#4E���l���J�
�(V)��5Ól��K]���$��_���;f���v(��`ӐgR)^Lt���$*6}N�E��Ք�㷥�07\����8���T��~N�߷�b�mo�B���xt��X�"��1�6k�(�U{�ɾVxy���e^�%w,����$+D
^I2�mv�8
U����:k��Z"s���WO:"�/w��QPVeYc��!'��r��hҐjA���e��BZ�l��с}TU��8�^�xWZD�(,�'3�d������~Wm�y�"�B�yLY�I&$��E�sq��>�Q\�V�����)����tv�X�:�q
��|�%rs���~"69B�{�e�]�,\��.L�t����h#г�m�̞�Q�e�x�Ĕ=9�N��`�J��O\���*v�7I��f[�]3u[XE����ep���	)�
V��6�~�����*�S���
���z��ŧ.�Dދ"��ڙ�h�9���ϙ��ө0���|��i�lڬ�����d�נ7��}��ލ�,s���7"#N=�u!`/�ܠ���=�O���n4-��O�4�,��!)�˵�O��}��Y(�@t����θ7�8��sb��,A�n7�d����Y��y�t:xH)>Z�
&B3���Ћ�U�,�=���R�M���A���_��*����ª��w�T�\�[䢪?H�4���PZpM�*��挱/�����l��E)�D�E�ͼ�I �Ib|�o`���z��e�-mm ��+�A����~�������G,�_i,I3H@�kp�c`���K��]��HJ-��yT��i� NH5G��ͥˎ�ʟE$�1?�VB�M�ܢ�,�4�׽ҙV(࢝]~��O�CY�em��\@�*<�oD��U��<h���g���|2���������~i�揤?6F�X홥L��9����pĀ.���lQ뭉A�¨-/C�D0:���g!ir[�|\<����a0�����V���ǚ�,��$���%���9N�)�'����c��B�(�f�i������Л����LDxf�2(6� Sܫ9B/�����ԋBԕ%�H4��	�t�J��9U
�//8���Uu_R|�~��<ۇ��%��I�\R@7���pӐs�-0#���o�e�#<��*�gP��#�r�=����X��
A�.���vaA��h�w����4���)��Sk�*4�`�;���BrIl�3��1��*�Gn�S���Q�f��~<���;������\l�����La+O�QM9���P�6�*��(��;�<J&�?���5�)�fHN����C�Y2N�t�.�K,ڜ_a	��l%�)D�DԘh�&k4^go��3�$sw�5P|	��o_1����b*i��9+i40"z(��� ��3 m��|Eh2w��j�g �~j�}�Db>GC����RB7���墦�'f�Vb��r�M��}�W����nR���%��xS(�jM�7�k6oCG��,1��մ%��a�6\����h4��C$}��N�%m���rO�A&Ȇ�aXM�'���Q�*�D��$u��S6�dp-��Q����i�$X$� L��X �����E��I����M���	�E �nQ���D|C�k��\���~חp@辛�E��,����#�c�36�.��m3Z�w�s4����${�cK��n4�2�1�;�O�oE#��ؿ��0I��������yf���8����߂RK�x�8J��_�@�g-޽���f�/���AwŠ3��y�dl6�T����T�b,iG�ٞ"H\[�o�rն��2�>� �/ug�	i�n1S��$;�No�8�{�y����W_D�F^9�M��OX��8���h�^�-0R�rN����љ���H3L-�8��(��%_4�◌)q	�����;��c#������W���}5=6{��WN��������:�3G\�{mh�H���O	����}�u<���o�T&Ӗ����7�9GMFI6ٿo8%���kSi��"j����@���7�Q
��&jY��O�y�#p��Ǒ���
Yuc����V�vУ�%��Z*�R�S��յmV�4�-/kP���^��m�7g|����i�G`�j��ǔ1P�s�wuv)g-���(9������l��'�H�5P��\NGI���ob�l��H�pO6NS�*4 ���t��Xh��ޝ�aA��/�T 6�Td�:��>a�I
fS�8�WYi$ 7T\I�W����r��9޿S���F��W�� P9���2x�,ç0�L�<���ʥ(�������{Xv���KtFdf)���U�����G7�@�{]����X8��6�/�Z�:��WEm�N{��5M�SgV�� cn<�TqQ�873=��l�'��b��q��q!XlxVHYEB    19fc     3f0�C8{�V �(y6�~h�Y�d{�41}��A��q4�=+���J+ȪТ�J~$X�4~ڲot!y��$sbs߿��˽
�9l҆[��9H�>��c<z~���1g��}e��>x����7$:���쉃JT��>�2j7�߁�u��;$�%�����q�nJ�&C�+2iD(��7sw>���e\O� �>N�6���(e����9X�5W!�}s����˩wD�m��׻/�Y��
���rxޮ�$�ɠH�ث���hG�]����wp�C# Zӟ��գ+'���ŰmSS�?�K߬.Y`9������G���(`z�K�[Z��x�+�����N�i���w�)3I�?�c��w����S�����"a=ŏ���NI�4'W����p5�<�EM\����1��n
j���H�o;�������/�̞I���{%��}u}[�";���k�(�^��Y@Oc�����Oڔ�4���х,ٺ[���U��ܑ�p"G�T�w!W�q�yz@��v�[��
����cWO,7��� ]�~)�}1�h�Q!�����$�F��Z���Hk�KG�h���Ō���_�����4n��"ꂈ�)?� 5]�ɛ���6��ۓ�������y�%�0�1Ѻ��l�<���[1�����&oV�w���xcq0��.�����r��X�f����m�u1Ѧ�V��&M,:+�>n���,"�Y��7"H��U�+6�w���.�	t�ir�ۂ��F���vns$%�9�]�S&�Hǣ����|����T������BC��d� ����3�~߷U�=)�+p��du�OG=�UbOb���YcNp��k�׼@�[�g���AW��
���n��^|��;�?	V�:��)3b��ZRJ�߶Ź�rUz�4VrBÂ+��6QN�ꦂA�3Kg"��; ���xQ\�Q:�Y*�٫U%/uy{�����S��d
W�R#�'Aҏz�.�;���b3�mV�S�