XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��a9��e��Yݖ����ʤF�#Ob�Hf
��p!j2`�5�^� �hη�Έ+�R�ݢ#�D>�FR�~k{b��GQ7�[�b!*WEP� �/g7�B�2p���i��c�L0-������d�h�I���i�׈�WB�P���њ��jH�t��y��h䦬�i�g�@�}n���CYL2�`{D������|���HN��jra��顪v[�]�k�~x8�����+���s֩�� ?z��ɐA%@�a���r��W^wj��P��aA�K���l�m~cB������vf��~�,�Gl��@�W-O3��iX��i���0c�ݖ>�Hkq����U�i�q�@s�
X̉��]6�9'��3��O��Ո�g9���'�2�cPẄ|��ʩT��\q��n��w	$*)�K
���JO��\���0��%���t��Mz��� �s��4ס�(�eLP��^�� y��ZfF��EpӅ���s�:ػ�ȿD
r.�L/'~�5���p��X�s3�I}��a|�E9���c}����S�JW1S�k�����D/�� �������k�u�Zb�?;�Ǵ�Y_z� A���\M���TG�,�'����Z�}k�&���Oc�]�`���n�P�"q0�N�a=�/�)���B?LD�L���IX����K����y�1<�=�fp�;��M�1sp}+>�~��	]7��Y����2�ﱬ�n���2a�2'2�d��
�ﵓ�&&�bџXlxVHYEB    fa00    2330U4V�%.�5��I�vUpo�=6��\��ƩB��G�2t��������{�RT��u	�0��<�l��G^j�d#���8�I;�w�n�\�$Lu��<��M
T��k��L`.�Ux�N�*�9��6tU�Mj���+r:�A�Y�y���pv[��TL�UF���} _\����YOZsPaV�Oi�Y�X�r7THZ��fhI��!�#��E�5�� ��*��@��c�R�<c4���1��@��ժ�dc���]���j����H�eq-t�z�
�e"~�F���n�����h�8�s�ojng�tM̈́�G�B���S��:�">H;�>��fX�3ߊr�T�"j�4|S��Mȴ��Xn
J�e�<t/�����TA�%ړ,��Jȵ�?� Ȁ��m�A��n^\v�wo�C�;|
)6>N�O �����_�ȷ��y��S��%#5�@뷨XA�,��R82�����:^��� h'Q�@����x����`�޷9}�$��#�Yn���C���՝�]��P��{)�i&�P�uO�!m�5����O`8����Sg�j�3[�*H�~��V��B
H*pV]�GPkϹ���w&��D�?r������#�hܵYVʿ�A�:��x��K2l%��F�'h���,�E�ԣ�����W�ԍ���	�Ys�ܤl��d�E�՛�@�#�e��5h�U-�uh��t�����N�9�Y�����̀�����P0��{��� �"E/���B��[�``�Ʉ�k�[�R�@�q)���;���F�@��˴���a�錡����t���eZH�2��ٝ��FM+ ��Tڈ��Gx�w�g�_�YB�P ��~\��Ϟ�����L��s��},ݭ�t���X�ʡpз�/J�|��G�g=�b��1|��|%�h}��2]h�$��kp?�"e���=�˘ٚ��CPr@� 3�~����������D/�F|�>����+>o#����q�qz���_RG�����G;���R��AI��$xy���:�p����v wK�����)��xL��Q�#���m+'Ğ�W�~����(Mx-�m�M�����M��i^�/�f
���^I�>l�v;p�	��?����q�m��� �s�ְ&s&�v^�1�e�7�D#�=c�x��6kEV�;SU��|�]�'�~�h]�E�7�gR2M���-�7��]��'r�l��0�0-˽���J
��9��<�ٝ�Y���L>�q��7��D��~l�����F>�>(C�t�.�b��t�lUj�Ž	��Gc�L��p�ǒ��^[&⊦���ݲµ8��5�'b!P}|27�b8���o��VuA��7ꈓ�}�}��{�����e9��h>vJ�W;�!t�(�C�������#�O7� �dAW+�՚ >>5g���V�au�_��t���AدE�v�Z��u�o�ܧ�Q?�����+��P�jp��E���k���Ś�R���]Íl�/
Z\�": z�m)	v��e���N.��S���&
�}@���]����8�*��
�J���f�)4~y������X�`F�jI Y���I�>��6a�@���Z�M�o�%=�q��Bp�Hi�hmX����]��3ӽ_ʌ��*�:r��rH�ԃ�k�f8��~�"c�@1��)Y!,C���umN5�Ï��@C��3Q�?�bJM~�A6�먈��p���Ȣ܈��B�x�ܙr��P������d�v%�-�P�I��W��P#�Ǡ�"'T��:������m��$ �s��m��V	�1�i���P�e�.!�<�a°ne~�$fK_#�Ӣ�B�s]@��b�[r����*��_�Z��f�������7$����/�WO�_#�#�����J�@��aɞXj%HK7,	%G�ń$�����G����r��/����x�\{��t۔1w/�Y��N�`	۟�J��od�)��dp����fp�`x;A���������SU��2Ǌ��!38��}V��])I����������)�_F��=��	���K �I[�508�P	U�X�^��(㊨�?���&�[
�s���Ŵ����o�T}�1H����3(
4��:��/?�VQ�S~|���aW��
\5����g\��j�����|y���g�f��n(�09'�g��f��Ï��H=��s�=?$�@6ўn,�4�Q����U$�޺-�5V&m�,������z��:�Rޣo����Wg����!�J!�7Z �b^����c�-�wo��d�щ���;BT1�8qb�Л?(�6[r���+�F�L�;=��HKߑ����4j�A��W9�!�gz��Z��ږ{�W'�u��|i� �(�c�f�@���7wT��Beo)gS!��}4��~���$3����S��6;z-\QD7�(Z��N����I��Bj�+���ɚF�$����;'Ҫ��3�������È�����{���%����l�t�xt�:�>I���
� f<���r�<Q���$K�/0c7u��2(�|���w*m��6�s�ҭ��l��~�����ܥ�����oS�܇}2�7�q����8^�%Za��?�űeԈ��ը���)p~��].�H!���<��;ֈ���"� %��Fg4sK}Kg~�?���C�aw�Ǯ���˶���Q��1���Vt�����M�SxuG�m�u��� �� �.*@9>���i�hL��u�,~�ρT��j'�#����y��8 �<�5[ߨ���,\���h�w_J��+*~����NQ���D��뒷��s-"��n"�3>�_b�����&_�;7�U�@��.�\�wP^��*:0Z���p���r��eiA�X�h�h�G�@��3��7�����l����&O����Z���Qm-��+�&tXGz��yQ������ _2|!�q���r�X�`��Hx�뿿%��N����Q!,2�īCO-:z��GxM}V�`���ΝvW�j��K���˚l.�d�Z��$P�MP�0�k��\���E��_ c}��K��fga}�V��>�m�ecȴ�fC-O���9K��6	^�y�mt�����;(��U�!--��q�w/sg/э�{��
�bd�2�X�8�k��_���$Y�*�h��\�V�R����Y��5{�F�/L��T�
S����V��t`���RL:��s�����\ZO��Q�z �ՠh5����9���4�Ӥ�]�J)QW�`���1������r��dgAz%��Gr\Te��=Mk���o��"����:�y��8���BI� �)�/&�oU����/z���(U �2MG~0S��gҊ�歠�ȃ�|	-J?-����*�h�D2�W�!�)�Ti�ÔN�ț�N,���-3`�4�Ṏ�)6j�6��wGM�:wvc�Y�0��.��|����"��8�RG�C��M�3�@�Е���8.�����Ѓ�n�Cs|SFO�BGW:`�����> ���Rd�V]Y޾�s#yw�;�x�h3;7�ŏ�%��� q�\���k��4!1)�WZ�����6�;����e^v������F-n+?X���2t���+��䓤�?*�%U]M0���:)�D�P,4��v�Ob^{�Ձ����y�eM��KC��B$'�(k���ye�l���O#�m"�5^�@�r�}% H�	�7��F��}��H]�Յ�y����2��`��5��{���Gj7M#�V��&?t����U��'q[� ��0����;xᲓ֭�W��	��@m.�KO����別��zه�ddR�'���	 �4a�R�|�}�}�L�pO�^�0�(�h0p]�$��im��a��T
F�5瑶(	�`��7?p�U�w�_���]����`�N���n�-էK+��4��R��m��/�~5?H��eǿI%Ï�rm'5��A:{�s^�?�pZ�7+J
B�b\ ��,�a��H�k�.G#����+�Z��b�Аv
�!&ڱɒڃ�����_��Epx���wJ������G���~DXpM!�%�����y�a��|ZE�BX�Ig�[(�#�hfcg��xtˠ���
��@�aD�y|a�A�˻�x�O���򂩁e���� �ر&�|`$3[7�5� �D�{aV���_�r�*	�\?�����W���^$�t��&3�a�VA�������;ml��_-��m2E�H��Yj�N
�iC�&S����%E�֥͂P{�/�|Uo)�<|��w�۳���0�S.�����i��J�}�5v�/��e���[���җ?Ȋ'N+Zh����Ȟx�4zZHƙ=�F�uA���d���8`���~�>��ո��S�AA�-�6��ڤ���]1�{/C��g� G�{a��\�X<K7�����_#(:��|��B#��f��}�,a��ٶ#2��j0�vFG��}�5��;-7 I����R��JJ����9��e;_�G2���l��滿�3F��剉)�"<����&`<��kn'��B�{�����M�*Md�r"��Y�z-AW�SJ^�
��^xG�o~��&���0��Y[J�O��՟&k�qO��v�%��7��a�:��|��իH(|�sE�� ����Kq.�&��\��|J�W$��g��&UU����T� ys�s@3��&���҄s�L��~_���71g��_r/]��/n��u�/0\���8��m�i'�Ik���E&����)����J����"�;c��b�3a؏}K��bթ8�2��	��!@n�_fg�8"(�������|�hĝk��lg`��@a�$T���z���hׁ�A���Tg+�X�f%^�A��7ԝii��1�c`,��]'�P�{J�`咐�1ؼ�v���E]��I��Վ����T<�)�O��w":�5�e��;��|����p�&��$�1����h�*Pv�+[]QT���1��� ����w�J<��\��C��c�LAɺ����/��D��Qv�Z�^@+����#C���	j���X�o�P�a�*�y���� �.r�ǣpo-����UVG�_��*B�T׈Y5�uO�0��q�����s�Q�O��0�a]/B�DZ�A�q�,1Efg���x�-/�eRYh���G�j����ђ������e�o��?�B�T5Y��-�S]WZD�1�-d3p�e��8��4�Ǆ��5��+[O]�Gֺ$qAx0п˛��JdAp�$>�C���H�eߢ�ښ���
���c�: �@ω&O^�����~�S���@��{ ���9qJBJ��4�%�X!V-Q?�q�:��Y�T����}�RC��e�
k}�F�T1�[*���U�)G2S�� �|�Ǚ@����s�s.G�~�\-�yY�T�=� I��Z���0`�� �ɾ���}����q,σ��UȘǒ�p�{��Ɇ��V����4)�M�x��u�2"1�]c�}�����hO�կʆ�5H������&�|`M�v�Q�� �'����U���,���?sXB�.�K�`��o���m��Y_�pL*b������fjU<w�A��g��ʾE���q�	��vx��Տ���3��:O̢��4�7E3J0$,ļ�z�9�}4�!��*��Ļ�hU1�N#�}[||�e��q�.F�S��i�m �Hي�`��ځf�Pe���a2PG;2�V�7�x|����h�e��\���B��cZ��@
��h�Ǣ����F�>�?���:�������'�)"Yd��D�� �B�R@��	���GPI����N!�����# �4�}�O%�õ�
����T����'h�!%/}��P����CL�ړk�(����Ayы�?�16^.��R�ba6�/�"���)�`���P1-{o"6߾�_�r'Hڜ�/��cT	�A0�l�P������f�S���4�dC�q��ַ�Eۯ�,��G̳y��{}L��&'C_��Be�R0V������,璖��PF�k�@����Hͻx�!�b��"�%�O%X{��rGe����A_f� ���҂����Z�!���Ħ���)��*}I��3��8�O�>���_�X6k�H��	�J4�6����i̌=ry6~��q��3-E��@i�U�L5����Cqި��6���$�Y���&\(�B�HԾ�>o�!ev�.�~�YU�k����Ǣ����꽹[)����|��~Qb`|Ⱥ���#�#��e�!i����:9l��@��޺�ǥ����S�|�~FZ�L�]h9sw���wsM�ӱ����6��L5O]�W�pP9��R�)�HB���M6�{O���1H@�F�qˤԬrAɆ' ��ƌ�+�����Om]��4��v���TP���e��ᯚ�Q�<��j˂�r�ٷtZ��>S��|�}H�S�,TbT�dђC��$$ǘ�r<���@�A1�B:6
�4����3,��@@6�S� ��HW�C�;k�E^�1F��e��Y'�<�u�&0&����wU
���Մ[�p��^�lV���	;'{�X�G��#� �����id����o�X�|ŭ�"�����@QRHMI�F0�>���S��������k��;[�;2�B��M����o<Uڻ�@��i�'��
,v���U�S,��G�@�$��r|'婗>E���b���'Ɔ�gL�2�`JT�CP�ג�e ���ڻ=��9\ǝ]ܫ*1p�Q�yH�L�j�0���O�CF�	t?�+q�O���j]�; �'�����f�qeli���on�JQ����#��u�zߎJ�'��X����۶e��s!	�A�9�{):aK���_��r�$��UB����O餎��F��*8*w�Qx�m:H��]>� _���̱��[!��UN�.q;�i�z<|����q���=����n�QJӐ��<&���1M�?���
������fٯ;�.�n.É�n��MG9!���\��5��=���O��x���p�#2I
��~ V�$���\�BϋF*Y� ��-��DT"[����)ZKz�ʒ=�ɌIPN�d���[��{s�s�����n]��Sת(���z6��Uj�&1���x�Ma;WG��"eH��s�<免4�`cG� ��ߢg���2�6���r3t���Mve��;(���2H~
l3n
B� ��J����=�H8��nX�sz������w=@a@o^ ~$N<���h��E�ν�1?�V�b��LO��xo�b���h�'�LU4�,ۿ.�]J�R��T�G���A�����0�����Ҍ��~]�Roc�Mj:X]�X��|k�Q*eo?w�ă�ڍ]OZ�f0r���� ������Bк]ƈ���U~ȭ�m�=��K�K���1�	5��3�avN2������&f�\!�5���jX��]_�2y�tZ�-8�[1x�Y��1�)8�=~B�԰��uT�[��ӏ\Wf����5��,��m�Q&�
�hI=0L��{�����h�I�﫱�2��]0�1ǋ�g�A��2�'�����~��Bj�(��Fu^�;Eۂ�cC+��m�ˤ�
;���+�������M&�<9�W��B�u��G{Tҫ��̆Z�
"v=]�F���Tw�Mɉ��i���Z>�{���{�E����m4�3_���
��\�ht������8|'\|�:���o�!z�����Rhm�lp/�k�&�EJ ��@Wk a�,��'9mc�?���΢}7��-�Xl*ЅNj�;�V���J�t���sb�I�P��N?�?���+��ۖj���W� +v�gQ�w��+�zˉ�^g_�*X����dH#�~�	!6s�s�ns�X�MV�w=A����,g�5^d���[��ן�y�n#�!�4���a^�o[Eml��|��)�xo��1\ֽs���G?l�ϧl��4�Z�Hoܑ�Ŷy
���)H]��ӱQ��t���Y��X�BWW�'7A^ L��.��V�"��l�T���z�r���*O�5�D��l�o^F�����l���E:W�8����B7M�=�L[ۨg]��lb�3�?���YZn&�t<r��W��8QF0�N`�l�Rp�y����c�A+@̤�u���h�ɳ��ՁESX�'�\��˾g,�U
LB�]C K�O6*�8���QS�m��k��� n�ܕeHV��\�@J#�t���
My���x�=	�P"ᵦ�{Y<��D�0��Gd����Sv]�
���O��̒fg��Nk��`��/�I��WU�q�'�6��w�og{��ǭh	����-`~�?^gW�0HN��uZ�����w� Ȅ����$����7���e�� �� :R�����rDˊ=�PZ
&�LP0���lR�9ngT�,+��/3����%�H;B����#�`Տ�w̢d ��R�z�t�d�x�7��Y
���_ct�t�A1��yh�@��ĽBݶ�ȹ"{�)R�	Py�p���_ƪWt�����B�0co�*s���}��#���)�+�A��	���АA�p_{W���`�'��H�t$	�[i~l�;��K��2��|/W73pq?��0*��5��������6�����x=-����BǏ���H�����j�Ap@����*�8��������_�"���g����GOqiM��U<�O2��2���22�������~[�<��E�_��b��Ϩ���7���Jf1)x��n>�a��¶�ER+��(t�V��S��3d�Z���8;�[�=�^�^�x93�N:TC���5�?̝�ǌ���!lP\8���Q���!�Џ��-_��4WXlxVHYEB    2175     710�ڎ���O��7L����0������-����| )HLDۍ�^[!'��"L6�Z`Ud+W�SR��w�P�,�o�'V�@N��d92�8�R:�zq��KЏ#�E#�T#�����X!M����c����C�e�����秵_��J�5��:�`:�zCq����F�\j�I��E?��史 �L�o��lߐka(Ҟs��(�P�R,+�����4d�z��� �`�z��R�M&ΐe�LV��i�@��GeQ�߳��s�R-���R3Dh��B4^g.�x�]o�"�
�1M��=��Z���tE�,z�pT8tyQ�
�Fs����}� ������{l��~lW/�O�1�?#��m!�z�?���_����?�ރ�tP�{�a��S�I�(Az9K?wf�W���D��ߴ 
��
�V9�(R�P�\(�A!�Y�T$����!D������?[<�6�G'VZ&��I��4�:��˖����%
��V��w�'J��[��������`0,j>ˋ��~��C9H$~t�i�)zg���3�>J-����V���X��`z!�m GX�]�t_��7�+v�%�>���K�h-�8��M��)�mM���^w�ݟ�,�<�e�	X��÷������N+�>���������H������O���
\�Im�(�Q�1i'Ma��:��\�=X����M��i������猟���{�緪�SN�m��u�G��Z!�&hyv�,]H7@*�\��J{bHN$�����E�[����{q�.��-M%� N�J��ʏ-�r��;�
G׽!�m��aXy��AZjBH(��<">h���dY�-T��o��J��+�"�t+!@���D�$2����D��DT*~���h�
������N�D���LM3�zI,l�#.���=��������쌣��t#�����.[��<�|���;������D.pV�)s�_P]F����o�*m��@X�G\?b���F|yug�%e.���?HQ�Lݞ��H�<*��vh�Y�<�֏Bg]h�np��Û1Q�{�� �����nM�A���5}��12k���c��o��6�+(7P&��u��R`���m߈M8v.Һ��"
����.(t�9p�\�6AG��1���A��`��M8�c�����`���Wp0���O�Fs�hD��x?�yh+���@��zD���r=�٩G+�E]o��\��/ҽ����y�R�Y��Ol*L��`���d9�1�9M����s�0}f�����_�����ߨiյn��K �f��Z��>jd�ﰳ�-�m�|���׼0s9ZAɍ׸D�w5v��Ѥ�Q�9�:��7ӓT���M߭�f�Se���n������ ��l��|(B7�UX��lb,��`mF}���}ҡt�:���A����)��%�Y�@��N��G@J��;2�}y�\O�\D晛���=�����{���EԾ/�	���j�jS��|�8͍r�'\7�w[HV�$T�Fh�R��$uKb馰)��\��֫�A�5w8Q~�جP}7\GT@ٿ8�^װ�/3�R�����wd�/��cQ��]���8}	��hH���/P�_'O�S����UX��$��
rvV��;GV��c�����dH���:K��a�{�ns����k#r�9B�#�lv�y���	K�����J<F3�B���C�Km0]�JE�q%d��k	)��P9�R�tJ���~26εL��E4���SI��io���h[�ˌ�SQ��°!eUO�_��q.S��|�I�