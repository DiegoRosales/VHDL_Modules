XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��O�u���]|�=o�oJS_
 ��� �(Р��Zx�|�$����P>���7� �:�Vd�?�2C��d Cr(�Տ���U �6���N��+��	��#��V��'8�QOL�3�(�7���,�!�6C�^ɋO���<�����M�~���R�p�E����������yQ�H�q��
z���p�M x��-���毉&�S���j���[�thR�Ć��Eg�Ǿ��7�N�Q�e˒��Hx���I�<�(���
�|���>�4�>\?@,1�T�؀Z'pz�3|�<Z�U�����R�T��#1s������/��6����:�E�gч?(���3�z)�ʍ��$y��ZT�����v����5)i��؄?W�cX�^���m�m�o�K��Y_�r���Jg�f7�YMǅ��_#�����W|L�.�vSM�<]R��� ���Op����a6�[�����/R�tuS�˼ $$����g5}&)���`'.�G���3S���\nc�_D���x�/����D0奢�?C���%��R�p�U��j�+=�S�YlH�&�4��6��*��_E�f�~`�>#�)�������gh�.Tm��Two�`����������\ԁ���gߤ��_MI��ZAy/��6����ޞ���Ӎ��8J�D��2�韻�$�~��2�ܢ!wP��uߛ�g���dF%Bi5�D=ΦQw�6�>����3��#���㮐�k��������<��`'!hP�#��f���XlxVHYEB    20d4     b00�Up~i���AphA�@���N��i��A���$ԩ=�o��^���4��|��1Y�K�)֘��S��H}w*�zؗK�ɖ�Y޶ D1�h��,�P��g�*�3�r����	ͭ*z��5�����иrH:Km�?Z��a��|Yr� �Y�>�.s�n����8j(c���1��=4C�e�]�}�T���_��L"���%�;���p�n�'�)W'��������S� �b ZgK���d�b�FR�f�C�i+	�^�u�(/׍k�{���[�G����4���(����ە,�Q[�4��2��x���T�K�Dz�7�J��G��� S>�
@�g4������E��������3����#��C"`&�'�n�FB�<� #�U�������'>ʁ�tP#�X��^�S����W�D��ٷ�����ձu�xH|��s���� �<�ᕥ=�{��>��� �Iw. �������7	����_����)�5�$�/t�C��2��5�:$�ܫ��X��)ˆ�n��� _��v��j>:B�@���p�����sE��rB�3*V�9,Q����"l1�M�w��{�<xzͼ7�)���H�E8���@d+�K�soKְ�n�|�Iq1$�� �e�Y�ͫ��r�Z�<��NJ֌:9!��? ���(ܹ[�UD�
{%g���
��͢1��m؞�gԔA]�4�9+H"F�2'��O��r`
9����Ԉ��$ hpˌϽ,*ò,)z'D�E�C"e\Ѳ�g�ĉ��0��H��Eˉ5���V��Y��;t�N�����'|#o6���ޚ=�e���me�/� ?��`ƒrn���ϟ.���bx��xp�3V�Ţv�6��t�;6���E=�A@/>�N;�$Ly��ԗ0d��U�<���?�
Ay���P/l��E���Y����l��ߍ��H�|	cЌ����s��@6�A��P��˫��S�&��F��!�+�����m��R5��wǟc��؍CS���{��]�܈��V��che[iZ��$v�>�#��{��[�\-�C�HǤGf��&Kdׂ*=��@����q����8�i
1�v�ţ>�o�
x�� ��6���$?�����di�e�+�ݿ(�Dj1�o��H��6!N��ǍK�\���F"��9��e�sj���0P`�e�y��I/�M�eW�_�n]�$�B��Q��D���?x�2�����H8��(���9l���3� �� 5���y*�ʵ���gs��l�pP��KU>˄���[9�e��>O�
K�8?S��ɻ*$��q���~�&^פX�'7q����h	V,� �	������ό�+^� Td�qZ�@�QC�~�f��}9�.��ŝ�٭v@���ץxO��X��ϊJ�?b��ud �%���y���^^V#��U��
����ƥ��E3o@
�ww�qغ��lq<�D�@��5�*���̿�����J�DĘ��Eul�6A�ox��3²���,c��̬�ְĦM*�Y���^t�T�*Z1�4�v�" �c��2}�6�C��s뗚�
$�v(t5C���R���L&WY/Z˯?����C�L��ᨛ@���t��ƃ�- R��Ã�Z�O��1�(.�QG��"ҟ�FjhR.i��K[����9.���T�w�O�?w2?�h_��+
|�U���&��y��wWa�Ɍ�Ͻ���� 2P�_��A��?=¯c��H��(	
�ۂ��h�V�.����x�V{�Ǚ�ML�x���<��A#gP�8vB ?��m��։ȓ�E�:ou�G{��N��}���c�^G "�}�FL�H*Z�R܇����t�F�F�$�C�WQ��T�*�K��P�E����a�QrJ=�����ъTղ�U&��ɿ�3���H��7v���F%}& z�%�mui4J>��v�F�$��	SQg6bGЇ��c�U�=4ϗd�H���RH���f��O]����<o�U߯��^l7���*�`Dʞ7�^h� nn��N�|�P�r;6u��G.�㻠�8��C`�
�g�w�+�j=^>xΏ�d�R�����r����8:��;R@���^7aL�9su�j�4ZTQ�K:������X9��
�ɍ�N�Z�d��v<u�}�? �O�����0�p��S�*�X�jD����yBS��
:�2�ڍc=\�� ���o���x��:�eqddպ��{�����7�'������Ka�-�=p�9N��n�H�˒V�	0g1s´OW˱7��P�O�s?n�93�c�ӵ�2T����0���b�l���ލFd�Ka����i�N�_�G	�	ٯg���e��+�S�B��c���XEA�������i4~5���{�Z����er磰	�<~��.k�0G�vҎ�j�!t�beu2��v�,�,�ރ}
��R����k����4r��̭I�8Ao��^ޞ�i�[�8o�����n�!xF�&�x]Iݾr�gh�=�\k��z��~_�2��ks8��v<��@�< oH�ݶ΋���5�~���0��o�M����i }	��Z�"���!��T]���XN����z��Ρ���Άӵ݊I�^��f"�h�@=��4���t��@��q��B��Z�80��';���>7i���5�>���2���W���4��$���9�KKz�$RMK��,�Н
tĴ�1_e*�,�x϶`��o5���: