XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��@b�\u�K-?_sYn7$�ι�ye$	ÿ8�%����u-�?8�;0!�
�ۜQ���k��d�����M2��I`��^��	ܰ�Úu�;%w%ͤ׷~B4-�.�'ckr7ʩ�ukȓ�x��f�.\Y�4�׀c�B�W��>I�v��U��]��ze����P���\>��-��5��h<DSu��z�C,QUB�������0��먰a�q⾘�&Z,Qw�Nr������4��r���	�|��<����`$&�!���ot��l��:�B��S����\Κ��KGr�3�eE�[J�t��؎����O�HL�U%��
j<�^�x��c�V����d?0Idb?f��	�[��6��@T�����c����'
��ƞ��Wԑt���g��tyQ�س)Q5�<Jp��Net��a2D�E-��|dxjMͫGZ*`�	ׯ�b�gd�F�AʥD�	J�V"���9	�h�@*۶�Z�;O7mI�<��x�����u�m 3B����Ȗ�ߖWM~�#�!`���Afջj���J�.S��b��9	r�����8�͊Up�U5�'�]���ڿ�FW�O�}�o�f
7���o���݂ܥjN�`^Će}6E�d���Z���Xw�L������.���S�K	��f�E%\]�L��C�%QO'�'�K�Ϧ!{iS�=�gLr�����L���?8�9[e�������Ö+������);�y�Y�R�����K��qG3��e���g��EI�{�XlxVHYEB    1835     920�7+�� �ec��{)��^��˕��|M���j{~���ش�(�}��@� ���T����m]r��R��-�mo�@������fE��iӜ��Ӕ[�ix��Ԝ�lTIMʃ[�ɍ�W�Kx���x|�J̣ظ�:u^58m[���ܽ������xX�N��O"��t`]�&���5s#M�LŽҩ�/}�Ot���B}����Q˙��]CJj�ϏB�ӈm��g�����q�Ү��m�Ȩӵ!*ƃZ ���A��^]L&��JM���K�����SdM�g�˩��,�E�|;�|:6�@�w�#��N�I�ɚ���,��b,��X�8��,��"�2l�'W����C
�������#�yq{h���6�خ��P��P��$�_\� IN�\PF	%���L�؃�Ҵ����q敝pl�NMV����-i8�D��<�웬FI6���s{�x��i�n�}��U6h��a�fnCD�#�E�b�{�R-!���L���W6��[�-�w�Nd(����q"��Dcwy��7[��!J������:.-F2&5���c��\�+��r+�:����y:!��Wf�c�z�crA�KV� ��@�s/����R^�Z�y��K�/��S� �p�Xp�[�P��F�(���\��ƅЄ��|l��P\Y�ޕF�t�����a�\�ƭ����c)�ܞ}��m{r߻͔��a�I	M�E�j?�+��4�h��I� |"~�@������bCفD���� ,J���>�����n�%�G�v�D��y�g�hF,��N�aY�$�r�Ժ�݂�7`튯h�hfP��Xp9���&�M/N�Y3�s\Db��Ae��D~il�T���D䀘�f1ﮐ{;$���H�f��RKC4u�O��F�����l����x�[�Gh�,^��v�2W��FN��?RzC*������L��
������S���C�MFy�u�!u���Ȅ�����k�hC���g3��k��%�
��BvH������>>��Eڇe��!�P��h���pzю���jj��Jc��`���@<�o�����|�^B��u�U�k�r�Y�ć���{��!'%q=ct�;��We��yL�&���غ����.������o�R�bQ�.������������a�e <�z�"��RCЫ`}���e����5�p��6��/�R(l@�<���v�Ph/���j0��d>���z��z�xM4̗%�F����1�@E������5�48ܠs��y���۾*ďzs����3�6�����+��Ko�
��Sb�
"w��Q����;@��GW�Q��`�8ش��7��pG���q�fZD:.t� 8M��&
&�[�}�lA���M��������Ӕ����fmFL���'꾡�s��w:A�3.{=�4�?H��Ĕ?n�`Ŀ���v :��e��GY���3B�����݆�0To�����_e�)��}yՅ�#�h���'��t��8s\B�b�>R,���CҴE-!xZu)3��t.ȑ{9�LYh��.��a<Ҁ��"}��sC���&�����湈Z:Af�N^増ε<M��aa���P	����8�`�F��Ή�h�7M2(f��s�S���R��:�XiA5BTڲ�.zD�*8<���^�����}���D�:��᜘|����jk.O�Lᕍ�#����\b�R�:������5L���|��9U���Q�=�9���P�i�7K���g.���XXR"�u��Q��}7��J��5,��ȁNk$�d� eC���j9.�����XK�ü��:�[X���fC�R��Z���^>���IK�^�E�{�Fc�Z��-�(�Y��Ǧ�_�KË�A0�G�(4��P�;�qƈ���8�K������g�5��*��c������q{��;�������dȍ.�H��S�6`���ݬ�!. ���BJC�)W���޼s��N�@��m���;���\NFJ}~>`��\l�=ZjAJ_ p��\E�xT� ΰ�95��->ʹ;7���M��銉���O�Bg.�i��v�>"Fo�	SըۓXOP&�l�e�AU����3v���PE�c��޴?��ߓ�ʑ����G��*r���m=�iG�������oE��؉�ĥt�2r+���A��Q�/�(�R&>�'�U����U�������Ǩ7=�΍߬�k�-$`A�m#^;�Z��W�gdq�}�<�2��w�l����ř:]�+}0��s�?l�5���S����#��=)I�a�Y������X�