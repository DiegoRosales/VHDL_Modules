XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���Hlΐ����D����a�o�.l����O|�Ȝ@9�K����`���'��D@�"��	,,`)}� d��D$'8���];~)=�u��t�_%w�]H`�����9��wF�E�����ɓ�s5�+>�vD��q�珉��������O}��P���}�w��3L��@�N������4%"�c!��?���\��>�FI8eR��Y/m�`������9&I��rG?��BD�$j(�#zڹ��J4�,2xt�<�|�,��=��i���b������}g@��_Z+<��L<�:�u�����jU$��z6���Q����dG�-5J���6�𸻎L��6�D�+Ds��U����΂�m��Q��mh��1,�C>��o���KT�p�D~��4��2},�U��Db���֌<�����鄕�s^�����|��Zァ�bM�k�h���Iu�)�EҤW�پ�0
w�%T��G��a�u;��ۚ�UM�c��.�`	�n��&� ���XC���f�BXaen����ojKt�5\Y<d�����mqΥ哯U����e��(�BN���n~�.��f�>ML��EV	s�;T�q�
�0Ap��ٌ�ꩼL��Cbm�V�!C�2S�#��mp����K���{�v�4�X�Y*s�P1��ˑY�,�Q2��[M�C8,�����I�E� �Mw.?�U�"��?��Q$^�����=�6�f����-�g�{��Jh���T
ʛ�`����rfnXH7XlxVHYEB    2dff     d40�ၖ�M쬊��D��r��`ř{�E��|�����S
��9�
��r��򷶼"uF�\�P�G��z���_��b�gj^>������+����硣6,qk�ӓ�\�t�:i�V)1�l���q,̰��V��	��M�G�l�-��R��|�\Z'%�05�&�
�?Of�$�pR�������Q�_���=U-�I���9��4�Meq���іvy�o`�g� Bg�#,8w�����P�K!�@y��b� c��>�w{d}���TvR:��Ep(zC`�m���Dz%�H�6�����n�^�ҳ����T��9�D�Ɓ��`���(�~��[b?H0����H*��N�x]Շ{�l�Vx8$6�M����X�,҅o!��P���Ԓ]��� ],e�^
�r�t�	{ƀ��|H1�������_:AɗY������\@Į��"������T�QZ�����Tƒ��u'��,��Ӫ�@3�������`���Y�v\������$:��fmk�a0XQt(oS4P
'##�Yo���;�3گ�+����@�i����(Ĝ��B�o�]ou��Zڢs�0���Ϛ���O�����X�����4Ө�>?���)�g݀HP�z�pC�O���3��tr�ٟ�A�tvb������̓2�f/۴�q�*I�B�8p���� �AF.����\��NJC��A�¥�ʕ�<鯺`u�ռ��	�s׆����P��W�=@����������������\
D� ��� �t��޲f,��e_ pFf�ξU��Z�Ih'����U^����f턯�u�Kd�"��cL�T�" ���c�&�w�w���j��{�jR��;�'�)��*P�̤D��M��M�/�e3QlX ���Jn}.&<� e�e9u���T����EP#j1�0:��S����!d����<�_!R�p:�)�\��������'�yӟ��e@�	M�>LCu��[��\I��x# .8��������~��^rr��^�����/1H�)���N3�����4D��a���RWЋ`�j5�W��w�E�[Q�E�k�a��"Ȓ{;=o������͂�n����5����4�ڳ���� �J�j	��$�#�Y�����9��xؒ���l��v��("�n(^�Ք��6Gm_����Ӯ*�%���8(ia��?� k]��z�d:=�+��KiT��Ǽ�;P
����֧�!Ѣ5��!�ֳ\���G
��
�X21U��Q+Ͼ���r��F�L��t������� ��ƌ���/�_C��}6���"���CZ���F ,���ve}�1�/t�
&��7!<J*�ڟ𢎠�#4%㹓�����G.Y/��vEG�0��H�G�v3,ҟ�_��ۺ�m��c�Gʑt�����{CS\��xv��OL��I
���R�>&��d�`*3�XE�J*8O6s9�Wo¤;({�\q�*,}>���:\+�U�������]�o�m����d�$������1ǯ,	C���
��
W]�ҽSL6���&�Nb���&gxٳ!{�_C�����PP&N�.kj5Aol"��&���~��\�xea�Z[f��m��|�9h���w\ǋ@��PCm{ة�g�
W�q��0cX����k���˳�i-g�ޭ�%�4�9��2��8�.�榴8���a/Q<Cw��4��>a�,��+^�ط�?������L�lW���"$}�vt<ZsS-���k"��_<W��LѤ��<��s��\�Z�����x�z�e@i�.��뱠�3@\��O�"/�2MKY������pК}��֙�����Y脖�7o���.�ZK
��
u��y�!����%�l+�"����_���v��&$��H�Qb6��	�@z;�:s��LNo#fX9ߌ��d$Q>�S�I������ҽ:�`K�wv<$��!�;��|������X�#��ɒxfW+��j��(N�X�p��i��d�ŧ^�
���򏑦M
�Εe9�]�߬��֯�h#� x4 d�P�6 �D-����5D�HBީ�g�#�H@X���
S�Ƒ@'��O�e���k�xqpFP��̟���z�wEД��O��)/'`�*g�evք�k��~^��n�0��OѽCf�l�.2@O�q�=P� �r,Z�A�Y%?v�2�$wϿ8�HmY-N���v�bi�a�����r�J������]Q����W��i����Y��ɼwAF.�h��<O�sJ�\��w��2�V�r)��7����wU�׆��m�����M->>ݗ1��*uv�Z	����	��oO�4R����E�}*Je�^��"�$X-k���a��{J.��.�FL�֦J�##m�3^z�q${�󶱉���o�T��C�A���UI�?~q0���O���^y�)]�� g��Ke�'Gӹ�6�����R��<������Z����|��\��Z��D����ɞ9�5��v�3G)��DI<%i��*D��F��lҔ�����Y��a�]����9ď�]�w�暪�2����Э�:�V!�-�|,��椴fɢ�F&�E��]ǵ��m�o>ҿŜl�����t%���gWz�
[�Yc�9*/�܂	�^<������o�B��z�U�R�zm�H�$oY�����(V���	�3�?zR�*���F)Jw^�f���m�C�#e.�Cʇ �2�\�!��4��Zi���������a��r=��z�>�NC0>%�Y��G�T8��P�:q�k��ce:H0�ć���f�󉉷��U�41#ȵ��v��O��m�9����v{��A.xCs�jpT�4�+3}��L���R����"����՝_�B"��r�*��v\3����P�nf�S�av��S�h��TWY���=>O'�_|��X�muP��	�Љ �A|�.F � ��p��d8.���Kv��k��'���5�*ivy��S�e��R9��7a�o��ywo�N�3i����wR I��[�Q��sL�4{�꧓XiJ?d'�q������3��3*E#:L�m	���]e^��}6^O3T�v@�Z�-߿����|�I�+�/y��&P^h�숯��	\����'���:��)�����[��ÚUe��}���U9��&�@p�߄eNa":�%�[�|�O؏d
}�c��=�V�k�I������1n�Dܐ�]%37W���[��G;�<��ۅ�H2);�e9x�;�_�4���;~!��I�ͩ��b��?GJ����Q~:��%�!E����h�>^��}�l��1���z��y�1�A�mrE�C�h��]�>(2Ч�;ψO�