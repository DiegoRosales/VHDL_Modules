XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��x��k3��p;&)�÷��B����'qj�?x��m�"]V:β�'�V�̆+"�~.�Τo
Xer6��_�*ͦpZpR�.��s?CL��&�S����x-I��xL�/��T+2|�ef�z�k6ɾ��B\)����yA��A����3Y!IA\�k��m"��4�<-�4yZk��^���L�ND�ɹ���s&�R���$���Cb��&ӿ�2��5� �񱣅�3��0Kr���
��Bh��N����M[N9��7r����#_��[�V^>�j� Vv�K��1��EԔ�`��گ~9 �f��H������YQ7V��A7��%~U���$������I���j���i����yu�o����x�|dFǯ�X���}���3$���w4���b̎��#���dW�W-s#[͆�aUU��z��?�*����)��v�MB#2�R�p]�c?d�-��M���^����1J��E�3xt-bz4�������!뺉��Y�LVO�1#���lN��M�dRl���ɍ�ɒ鏿�ό,/��oWg�v�C,$��y���4w�l�*�G(m��M�+�P���������)�<�,J?��:S�$Ou^8;b8mR��ƍݶ�TE��|e-l_�`�:�$1<��w��o�;�[�?d'��)��`��f�*TT������f��}i&�ǇV��ΪD�/r�-GOȿl��E�O��>�nU|�r�����&��X�2��tXlxVHYEB    18c0     850zkvUo�����F�d�����k����"��f;y4q8;��Ʒ��Z�V�K�]RF a���v�9��?`�>��t؅N�AJ����윮�������^��5�WE��w���Q��&���#0���ƨ%�/:@7�#$�C2iP�>���J��;�D�����lq>�Ri���3��؉�Zן�%`/`�����V�1�� ��#ӝ8,C>�5�|6�-�	�'n	$�zd��Q�+&Fh ���n������6Gz����x���R.^?��PJZ�6��i][��Mn�u��6C3�	��_A"�fe�P��f��_9)v��o�͘�:Y� ��{\
��r�����:������^�>����d{���
}qm�/B�m0�V�,dkBI�Y�=0G�4/�;��Մha\�5���#~2�N|&xz�k��k�Ǔk<�Ho\^"��Y��w���\m�a�-���O�}gW����D���;���9�)�3�Ճ�����;�/�N�iE��o�eM���As��y.$]�.�#��ΟzB/S��#q�ٳ��(�(Qr���[䌸lk+�)c��^��.%D����O}̸�f
ܛҫf�J)�m��q��ӌ��~mA���W�G*�Ȇk�,R�1
���J��"u;�Y�H֩�a����r�ƬN�O��'t��]���#��h�'��?6Б1s�. U�!ei�4_/�N9��xD�Ox�.|�F�Jek�Ȍ�dȏm�ɵ��L!^ý#A��E�eF�SRE�|�?���.J��Esv��Nң���NM������;�E�kt��k�4���v"���:�4R��*���$aB"2\X�n8B&G�������~]ƽA��~T$!,iwT669d{����7��atX@,�񿎸3W����;,(�ף싙��*k��P�?��� N�/s������d,��B�}�Prӳ�N��e�T�M� d�R�:3���T���%Q��?e�`>s��)�%+�v�N1uO$n���9�Y�t$c�V=��D��zC�b�sg��Q��U����3�+
.i�JZ�ʔ���5�ɞm��ҝ�سhڕh��}�~�o(A�Xsm��qF"v�8����{� ?άT<`k�(&k�u=��5�#�����w�'�ڑ��~�@	C�6)�@'>�ц�.�g��@P��U8r3�Ē@�X�̘{7* �_ס�X��ΐ(�)�}���*��U�@������^�h/�]�-�q��'��"n����u��+�,����ekyP+B��$ם�vpA�J҆&I��/�l5�i�����MN�J�/ڹ�ֺ�ǲh�*'�HA:�Z7�	x�*�F��Kڷ�	qw5"�(sX�*���]:q�1)9km�R2E\�|Y��?@e��G|�T�6Xm��n.w�:-��)Z�W��8m$z���VX��R�E��k����&~�~[���b��q�t_3O��	����y�~nf)��4R�I���b6nަt.
�#f�i�ԡ��WpZw�Ďtd,�����"áp��x�d�0���t�}j�r��rW��b[.Z�uua��oW��ɾY�'۟w���]�z�A�X�y��*�k�s��`9�k�o\6vqQ���-v����"��E?�i�7�P�P�ӄiȣ�F]Q���_Jc*À��Fq�(7C�T�1}4FV�8!E��?y������Q	JJv5j���9�V����9���ë4��k����\`��E"��(�il���M�l����u?����zI���D����H�rSI���F��(��6��۸k��$~��5�Em�s�1?w_OS�tiY�XI����øś�L���]ә��h���I�0���!R��~=襏����Í�뎊ۥa�*�?ms��e���s�X�u@d��z�B&�-�1�}$��2��[�H%��� -��w<SU�s_�+�sbCqz��F��y∛����8@�X� �:W.������
D��\QZ���y�;F��1B�MU�]M**"�A7�z�LK�7�
�߁�n�w0��k�*y���;�EW ����.���掐W
��҄���q���F)��o`T�E<E#8�1�