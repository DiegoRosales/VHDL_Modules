XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��p�^�6� ���-��3�{!O:�ȣ8�;�|� ���ݽ(HFs�uky hZ�Ӹ���H9���(]"��{���H`�����kK�7̄/�_!��k�VEG������G�P@���mc/��3K�_�cz�lc��̼���?�T/���hA�����E��e)��VVW��{`	f��e��4Q�'r��8��"o�y�a��)�+ұ�	���NR��ҫ�urWJ�,����@J�V�\.���\P�,"���֣�U�G�Y�;�P�W1󩏙b�1��Ӎ+;�OǢ6�5�m�k]����uq* ?���R�-�a	<nB����B~�B�K�b9��}��`�P"�"c�,��dz�.�6�r�����@]�k/���`K�h夀�r<�"̆��%��;���o�S�����3D<=�N=L�R�[A]�������'��d���f΀���c�(����攆G���&hJ�[����:굟��G��B�*�eod�u�v����,]��aF.g�I)�O����M(}{� ��'q�x�����>�����Ҙ�^�&�ևa~=�;�:�t��,;�v���)[$�I(UL�Y��^��>Zv��z�5����ۜ���d���l�je������L�z����_�"vU�����s���Sh�^pAv|λ��b����_|;�3��z���X���L�;������xkU� Λ>Wv��
b� ;�B�w��hC��˪,�SK���� ��/��)]�t�XlxVHYEB    32ec     940��_# BWl �D���+��8���s[�O���(�l���)�&YS/r`�!��f�+�ؚ�]���
T�9��5���cwn�y�/�Y��m�g�]�]x���d���K�� �g��{��!��p#&K�c��>Y^!|�{�e6�`�t�`����Ja�����R���Du�Ʒ��#D��Lz}BT����ׁ"�R(bX�&TXd��GTs�\�pi�/&����6�W˝��֦x�ɕ�������یת�����O���1���<�H�r/�:F��SH�q������+ ��
�̀P��߼��Q\�T4`g$�B�`��A��F�tNpͪZg(F��K��-�hn�a���z?V���m�@)�r	Քka�ͥR��Wה����� ��ZA��u�܎p��U�l��M�`u���O�*��*�k��|5��ԑ�X���Z��1����pu��8�m����C�.��e�@��"��+N�M���'��J�sڔN�T�ĕk�Hr�Yȿ���/�I
��4v���5jij��X�d�[4���]�o�s=4��1w���dV`�RlvI^�~�h���2DA��&r�c������D���c˷�"O��}�C3
�H2�j�Q�{P+s�ol��}�k罆%�Ӫs���e�h��zS���K�Q��S�/f-;�~l2����aL���0b�pJUW@��n�]H��1���@�z��ν�NzzV�4o�O1�ps�i`����<7��s�l�*#@Z����^D,�]d<t,@'���XX4ȮgAU�L�l|��-�͠H� \����d��H������h�:ú��}�7��������^ԅ����T�G����`�r�T�r�����w��R:�zR�IW9��{�C{�,{A@]ǳ)�9w�K&Xސކ6�v5a�K�RZU'$%����s��\��{DH��Q���I�"��f0��h w1��ס'���%{���ܕ��7��~�6�n�K
���۔���>d"�8v�#L��}�Y�⺈S�k[�w�J7�.���c�X����J�p2tRdGi��3ݜ@����l�#y��Vmo0zd>}?�;�ڳz�E](�ڲH�}}�t�H��y*�[�x�dmG����s��q7�z��D�;R���5��8�mD]`�Ͼ����$�jdR�o��&P����B/�� H�y��8A!©Ȼ�$xI���0bG�֏�2!�T&�$8;��}��]�GG6�>c���>@L�Rk[?Ʈ�i��x���d����|&5ѕ]��Tv���|��lxZ�䗕���/��ѠV��:�����b=��:�����`��sz��ZJ[WJ���tȸ�Jl�QQ���	d�{Ԙ��� �T�b�7�B��}�Sa��5���x��B	؝K����B����pO�}T�Ù�~1���N��Tzƾ�u]\D��{�8������tBe>�S<=~oH"=�v�����o��m����8�͝E}R�w�K����&�Q2U��7����0O.��,L���ҢN�씒
�st�Pz /�="aV�.,�16v[���p��Ԇ��?��U�Te\�J0���&�5s|/˭t�ԧ!�WR4<�k@1���p(8�m���s�~Ƶu>:�#�\i.{���ȫ��7�;@%���������>��J`��G�6�Ի�!Ea�3M��J�]ص���ɫ��FH�BI>ə�7N(^_��Ŧp��|�y�菗��z4��KZ
���T������H���j<NPs�9�_\�Id�KI��,��O&	�� 1�_���VX�0s�z�����č߀�B*>XgA0��~��#�%�H�Ş�2ooc�(���.@�ྒྷx��2y�ޡJ7d�kd��6�+���i&�g��G��t�=�v�/5�������������a�.�)��ږA]��Egk�27�VL�]sZ�5Ol�5W���+&<J�Q�L����h�x�l6�Aۙ��oŖx�]8�^��R���m-�V�0 w0L1`A�y���'���X��� `|�0���^Q7em��!-)����]�OmTyR�x���!�֫���5�
kg���ŧܙ�1\".�r�Ԧ��*,��}`a�0D��TÏN[o*I;��њN������:T���4�	�_�.`w7�t�-��C�����|�P&�#�)��S��K�X��BN���1#o��f�E�u"�-w^-��@�A8�i�+5�'�2��d?ϛ�ghZ�18��%ٰ<��#�<�Bgʇ�!���:�o�Q�Pp�;˵�]B�:ZU��Oj�6Qޒ���3'U�YӴ��؏�c� 