XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����i��2E�ᗦ+�s�O�EQʋ[�ru�׎��p�T�$/Szx�X�I���4�)\�N���[��\�Sw$&P�Y� ���&��]�Ex�dr���8{�_R���Yc�8��A(��0:�����m�"��Z �zѓm�_�t��:��f���j-7����o�U�'"�.K���d�W?Į��f�D����+��ymZ��E�p¾�/p�B@~l��y$���h���J���o��M��-��|p���r_^5Bl�uՋ6[NB�V@�g�Nygc�#S��ѦҲ�/��	��9.`d"����a*�.�*/�hN�K�D�з
sFXrN!�9����m"j�;XS�h���2]�f�A�,��z!�ű��|ʆ�K�s���$l�{��~��;>�Qs�P��~*�<)Ol�"�C�+��Ų��O �]zB	$]Zd��[Aw��/�@.�
�l~�ݲ/�۴v7��싛�y�5s�iӢL��9n�� q<�,07c%\�.�R�{�⭠m��5�W	��^�C���r��>���jyl��uF*��a��|E�.W���X�*b�ց`9���c���(�`�����`���#�	��p����p䱤>�B��+�d�Q��&�bL��B�����0A\��  Cs���\{��}�2�b1�*���û
L�$��x��Kal��vW�ä�D���aDo]Ă���B��]�d������u
�1�e�J�#���c�x�L��L�K�����]о��XlxVHYEB    2031     b10�`׉��*ϕ�@�^{k��4S�������g�.�F�Rk-������7�n/]O8�i51�G�roRFWM��T�Ey��45h������!HBe��!S��0���w+�:pz3�äi�c�&��d
_�l;�h괸��8���*܆��XܨǤ�GJJ�!�]��dU�L9_֣O��s�s�"/-�����ҞꐽA6�Py��?���r��[�j68�C�ϱ^����/��<_�Ӭ�Uk�O��(�G�J7@_z�h�g���u��p��4u7��H,���@l,}�H���פm��i�to�Z���U�F�e��)Z%<hvʃ|�9��+s�O��&N6�:����CD�s�����t�Ó���d�m��E�����:�=��%��x����crk��r+Y]��%�F�6(&d��k-�Ɔ|�'g��͌���]���6:�n	��{�����M����G��]�銪7���&PE��Ԩ�&�\��U|�+̫�f!u%'��'���Lp����N]���7xP���>� #��7ͽ��g��+x���q��}����w}±Ub��`���d.���2,���qk�T��KB7��X>o���#0�y�|�Dۨ�#� ��h��}Z��恉�͈�@�n@�+�ҙ|ARK}ݣL�r�%e�$n�s�z �J��2�d :}G̅�sP�5P6Owҙ��q��C��M�s���q(ivI�ϟ�E��q`�&I�kN�O�Uˍ iNZ=�0�bm� �ԓ�]w���~+�H����Y�X�[�Ki�Ұ��m���K�hAxD�`��v\nҷ�1<@��sE�R�Q��6ŦGi�El	^ۻ���8�3�=aS�e��,N�i���NԷĝ	�0zV�s4:��l��4���;5�,�~��]� W�g���p�\�^i�>��V�>^��-�B�H��?cϋQ���/+�>�}�3��?�W#��Wpї�6�Y�Gy������W��@Q�a(�LN��k)Ǵ7�W�.B	���#i��O	pȢ�[��, "oU �CxdDQ"��g�Hij�K�Ӛ*�tWr�N=�7�D����~v�j�C�[�N�,��5��^6��VJ���:k��Ot$��(�\Dc��t�ӪR3%;e� �y	\(�v��0�c�q��~���K>�d!�n,y�j�$���������~@�Mw��{%����S�v�D�|����t���R�c�J�*ܛ�YUә���1��m)Z1�>�E�\j����>8�;3��)i�@+M�5�C��^���$AH���l�x�\׷�X�>��M��H}e��� ��
x�Et���4ʊ�!�d������ץn�:���m+��c�ȗ�-*� X(9��1n����b���0�����C�m*GT��-2;��V[F`)�36��u�!=%�ɪ�{�()%��_}F5C��7�d�=Km��xiÂќ´M	�jtM�"�|s�9�۰��g�X�V��W�y�N��#J���5�� �~��B�uJ��vj;�F#�pkF��2¨^o�֜��2!zHD.���n�/릓��ЊF����i��y����&3��/Z�ۻ�h-r!��EO���a��fe2H�9Hb�������=�?z�|W���l�C�Q1; �M�Q��ozj�N&<ta;O�d���q0��{�q����Gs�=�����EH��0HN��N΢,d +J����ukY�t0�^�F4��id���U���(ȗ)��[&�I�^Ğ��2Ʋ��7�k�±1��R�ܔ�A2y��?טG|���B�b�s�Z�a�έ�(|4M�`V�r��up.��T��y�!��X����W��QYnM��V�zBYS�1�[~j�kC���,d�7���*��f,��Ť�]��pb[�7&:q�	'��`�	̿����_c����S�*���_|��6��	K �m�f ��)���f����\L��1_�̧��"�J=x�>T�l/���;BT�Zhj6n�G5l�)�^]=B�Aah�ݱ�t��Zf�}.�%3�����Þ����>�2�Z�G'�wg�'+"^��lr��W��O���ߤ��c�o�6�:`��K�mz��:!�9�..�3W!��,.��&�Y��b��,��◛��o�53���,4����MʈyKX�熦�ͮ�&��x�īO���J����"��	Ն���^�4Cs�\��zU2Vs�"
���������֦2��Ŧ��#����I�.r7��ʐ3'��}˰��/�#�����5�]ǡ)�h����1�#Kin�y>�Qk�¹�D9P|�����l.U���M�j�	@�>��Y���
��b�6��_`p�����Bv�ҞUן[cÁ5��Y�(�v�ng�Fxa@"�)3��_�FN����?��a�nF�_�d�^�k��Jv�t�(4���
��Dx0��@CjC��@�ȱ���hL�:���B5?� �W5;H�	�����|��%��� ���c�|_	�sA�!��I-)�'V/�k�ng��ؓ��ʛ�&��EN����6R+ڂ�}�|!�.��}�a�r����6-FcA�rb���o���'!#cr��hu�������O�x��vT�5���-�m�MT�K2QHõ67��i��FZ(3�T�$�ݨ2��蟹 ��K}�8���Vp$���Q�*��B�'~�:���!�=��
|
����;{�̼+a ĲS��!�[el�.Vi�G��;c���ir.��.���`f����`y�[�U�
O�G����-%-���T�԰\]#����?����	����