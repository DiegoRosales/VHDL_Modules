XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��I	�(
�6�4Lt�Z$��z�1Gz�~{q�ϭչH����|w�x������+�~���˭R�C�d]�7{~,�ـu�a� ���$+��?�y�6��V��}�x-H�7n��_vi=sEy�3�Uxk����	������dG�t�����W��t����)&�r"`c���l�4���!��	��Æ����0�D��޽\?��Dn��Ds�+����D� �G`w/=~��Pt�Y:�,N<�"��NL�M�F ��bڬ�nz%�}C�';�s/���'(�� ��,�eL������9�j0� g����{ge�|Î&Y܌)�Kh �Y�������e
�j�Kŵ�[��}r�X_���W[Kp��)���
lM�\�A6�z���j�7	�*�Z�e�t���Z��D�k�ec*�"�d����Rx�����8I�a��n8���F�f0����X��L�Fڪ=r���M+R����P��;�(�⯰s�x!aK&��t�������DȂ���f���"Dl�L�Y%�b=%E�Ʊ��W�<]�f/)"�*DM;�F�MGb�G~E.+e*����\�`M\(ඒbt���qA%����5X�ϕR�C���7a�p	���*������i�>i��_|ΤS)��Q��Oڟ�I���pZ(���jmg:��O!pEǻ�ji��G|�r�*8�B≐�^�Uy�� �s)t����a�[$��9�K'2���q7��H�_Q�kb;�4s���r�|�9��;�-�dXlxVHYEB    8349    1980@B�/�g����p-�7�Pyp~�X������.	v.��_�Ezm����O�hl�W�#`O�= z���Q�=@�H��-�o��a�h�:~�`���=��SILv�*u�6�*^�������{�g��ӭ����4"F�K(��1��P��=V��U\���Iآ�W��"�Vq�/�/@%z��ok�~R"�@�c�~�2�������l�mf�
邏<��ع�Y
P���zn��氇'Y~�]`~��ӽ��
2���P�0j����Iɂ� �\�N5�h����V
�gy)�0�z /L��A��Ԏ#}�fq.��IW��z�	V� ]�'��ƍ�����P��,���_TS&^�k/��>�|�'#T��_G��?�˞k��]���������7��h%��}[4V��5�p��+����s� �K�黢�ʄ̒+"�Yj�2��|cZa�����,l�Nl�I�����'�?�>K�	���g�xF��Hc��]���?����-�b�JT����i1`�W�/3�8�!T:Q?ż>s:jȆK@��W��5*�	钃'M���I��<�=_���Biŷ���XQ�b^@�p1��H:��s��T^*�ο�� W�r6+�O�h�#�?��d	a�#Ц���>ђY�ÄCS�>�gZ ��� ^|-Z3��|Ӣ�� sFC3ڧDv����^;�M)�6�V��U7�1�r��4Q�e��^)sD�cꨰ>]+6cޓ�~y�1���ˤ�8����h�U�|C{N=C�D�]�E!^:א�o�J�_I��DxQ8�,t��Ș�v����}VIq '�Tb�1��hz4EJ��p.ί;&�<nK5;U���zҔ/�u�Qe����P�����e��^u���,ռx@;��aR+>,s��N4�xSl� x�Zӥ �,⡸��CP�0`�!.|��	�ߴ�������
Sn�N27�()��(nmg���	:K���L���9UGRm��6;�%=��z���M�,>$���u{�|�V��ڏ���	�Q��-bUE�&���>7��C'�IA������9���e��q�7oe%M[pm0c�8#`�@�n.P���Y8@�ށC���2���E�3x�qB �l@�'�p�T��K�FGԁ�%yWa�/�} ���o�l��N��nwN�v��o�j�R�0�����',=�2!'��c��Ϥ�=q(\��Z��4U�&�$D�UN����D��r����c��B�B�J�_��j|^wO�]�T-��c�VS�-�'?]��Z@ p�ڭb��G�7BT����G�� %�k�'�g쇲7���� qXe*��8��lT�M��I�ϟb�� �ú�Xl�_b����j����F�o����ې�"���i�=�=R��l)��`u��$��O�k;�kԮu����3�z��Okŉ1 E�Q�� ���h�����\S�(��ʢ1�^	3���f�}�kN�͏�P$hj�Q~Uw�_^�k�����T��	���]2�������R����W�қ�E�+��G��)��W'��]?c�m�68��
v<�)�B���N+�(=��ɬIL�f�Hr6��qG�l��;���yH��K�)��%O9�$��V��g��)�*�*C(�W���%}3�|k����)o��4�^�ފ�ߚ2�}-Ja����2ޔ''��F���Q�`�a;��l��,��<ݩ�d6Z�L�ǃ��n����%6�e��'�3=�zt�X!A��|f�h��8���{tZ;��-�!$�О���|��=�<P܃S�fe��$�X�x��4�>`�ċ~���S*!$� ��;s����=����?���E��0�".F�ܓH91~V�#�]4?w���P��50��7"k�K�s|LFJ#��]���0�b���G����ow�Nw��!|�=�ϻǐ��n�#�YIv��UL��ڭJF���x���#f;��7��<nw�$	ƒ�%�����hu8c�R/�i�`ʙ��)ǒJ@�T�=��.�ߋ�4���<[~ �kx�A�）��Ћ\9kq�����Δ�:}>p�9�8;������R�u���Ϻ^<�y����'|bR'n�(�
���΀c�UkC����ف���A0�?��ͮ��@�Z�We�U��*�N.�єX&�mu1o��"��U��(ab�Օ:=��>�UJ���-4.#D��$`LL��jLɋ5��,\��O� s�+x8L��C�n��B��b#�ϣZ�axM�*ů�P�O�I��ǰ�Nh5 {�v��	��,Ng(]����ԨQ����vo)�@�>[p�ٷi,ƭ:��%Ge6i4I�����Ǿ�4֟;�9��9�oyT(w�Ŕ��+'}Y�N��gԼ�.��&o���xN�6`Ie�ua��S��>����+N�F_�����c��wg�� ¾x��x��I�%\�0C5� �/%�i&�!vu+B�
�2]2����M�iR�*��M��[ԋ��1�t�+;��t|"BY�z���Z�ã�@[�[y�*�)V���D�K�M�'uA��v�9h%U 	�q��N�&^�|��]���Ji��u0��s	6ڄ,A��q��L>�T=+�-���a�ڿ� �B���	���|��PrL�)W��u:��%u��r�\9A����<�)����T�.��i�����^�xv;�� �u��ĺ?�츜��
�"�x�,���e�o��!�N4@	�\)s~Q G:�Z �����H�4j��}GgHnʾ6n�@���K��+-��T���v=\�hZ�y �E[I7�[�*��\�q���㲧�*� �6����W���))�c<�g:4��|��9�=�W��z%û}��zg;��%�M�vvHY�\��v�1a�o���(8�y빷ϗdC��f�L�O�&������0ð:��d���/�P�<�p@06sy���9�K3V��=�*��6�4���`�t9�s���}���*Y�E���?!�4)aѷm�4cwF���1jJ2b���ReEh��|�����vb���o�g�՛\-}�z�� �i�1+�^�=���0>���-=��a��������@8.���c+�����A^!%�.�,�Z����l*�{M��Af�v��6�g�ښΕ���C��|a��N&Q8~�׍@xZʨ'��@"*mHX���Q�:(�0D�Wy��law��u�@%��J�����K�Ҽׅ<�K@P"��X���oyuY,]�f�`�%^�1���M�݄ ���W��}xQ��$]�Jü�%���o��C_F��,�10��ӂZ�р��S��^�D����%�Y�GV��!&y0��s<ɢ�UNH+Pc!h:�����+�'�'$�;����|g������B����ui;Cq�vgp�t4Y�K:�?g��C[���Z��T\n�K�f�}����7��x�\�Й��R☱�@r,�H����KP�JT�E>s���d���<���[hʊ;d�x�n7��������8��#�MY��9ɭz$v0&΁��W�	B��>�;^��)G4Д�&���w��$�pT�ϒ�,�Q�D��5]OP�+�S��0�=h~zE���L :� �^P�.�����]}���.u�����'��[b�1�=f9�Ѿ���eỌb�5�@�9�'3b!zY�U4 �#ؑ���:�R>��?n���Q����C�~=��<�8c�R-��v��YU�w�O���-�',[UnL�:�ڲ���1Ղ�@HO�A���b �8�C>������ѩ���-��X.�ʡ��g�D	���X���Z�u�cjnyc�+I��U��Ò���B�mgB|���2qR��{H�si�&_�^�%��#zї��W��Ta������aG��F�yDݱ�9�*+�ߏ4v�Y��s�k�(���"���p�E��j�I���.�ln��u1&tٌ�z��,�Ѽ�-�q�ꇈ��b�&��
�,L/�o(�R	�m|"��\���� ��N��t4ee�!�"Z�����A?��5"c�Y7~�[/4��g��I#%3P���M�1^1�ts��	,�=Lh-�m�&�,QkN&|� g�¹���D�����[8G9�r�A�C����-�����}V�_��d�9�a3�(�w�Й�~�Pw����E���#
6�XU���;��v	�B�U�R���"'U198�K��mաR$z��@�3�?�rV_�R�rT~˼�Ȧ*��F�Ki��B5�G������b�ծM���+y#O4� u�KF'��WA�����"��H>����d��m�̥��z���I�Ez=g:e6�_�C-��|�;���]r|�[ĚdAKkW�b���1�ˤ�A��	�՗zH�-Qi�vj	b�����ɼd>*JʬY3�6V-�d��Ff�he��r�S�A�_�ʺ������1Zl �[�A��U3�q>���\�A&\*b��QZ����P�����W��&z���������C)~�@��:����ny�Vn?�����I���1Y>݁�o��J���F��� C���(DA��Qr��������՞1��}o�2��<t1��>�n���=�@TB�"���}P�^#�-[�x�̮v��;uCh������Fna�t�(W}Û�|���ms��<d��I(>�~˿��$��_Yoa��	�C�W_c\>E�;����6^#9�q�fτ�Bb�kMB,���ݧl���QU�����c�]U���{c!#v�$5=��k������e�fpu���N��{��[D/F���O�N�'�d�r�:�Mbq�v�pW>����<����ÝN+3���K�:-B:m�����&Ƃ[���� q�b	�.t1�/K��S�Q^b����B�%�1�7�$(��%p!��P���z���H�[�.`,�~;/�'���q��[�|X9�ğ��ʋ ^
�gv��eQ{��<̘�,ߟ�#�뀔^'�$q^ڱ[G2��pEc���p�NM+��6�0�U���1w�tX�9>�����"B�ٚ���L��H	Ȏe�C{�$Ig�'�W|LC�:��������H���a�#�#�W�4�8U��<v�l6?Q#�ބ�I��"N�5�ʜ�`U��Hqo���:	3>���W���jg
7��j}���>�Gw4z�>��ʳ�C���MYf̓e�?�|Rؕ�  C�f3V1I]��:Xs*
����Z�#qI��{g����n����xk�x"I�&(M3�M����
����{",L�L������4��If|X�&��'B���B�<i�"��)?�QM��-1�Vfq-&IÍ�z��l����-��1۠�5c�7�bY��F�x�q�O]��3�5D�p}
��XK�q���	�R�4� b��h �>a"g�Ex&�x�Z�n��Nv��{m�C���hBX�$M'5=C�F?B(�2�`�u����+�Ft�[��SPɨO�[ל%/�G��A		�Y������̂�WiQ�OAt����"{�C��!�O�^9�ɸ#RJ�.�<�/�G�9+��H�r�c�l��׳X=�D/me?�A����K�1��e�r�� )��
�Ȋ���;g�du�C���������5k�-�4�N�v�҇�]==l}3<a~S���1��+}(�� �.�ϴD��K-*A�\I�؈h�6��U��bT�����,�/�^��<���n�Q{�I�<i&:r����x&�>9�K<�ytId4���eWy�z�T��5r������uȨ���j�^�g4:M����!�ݮ8�'�����ݚ2�Sͪb\R�h;�4K�;�ya�����D�G��Qݟ��\��V�M:ls��Qxo�CF�	0Y-�E[f�����u��h틚0cB-a6w?�ֹ�2Û�� ��f��
E��g���c@Oy�3F�6��؎�ͷE<�=jX���.ږ��жCbo�/{����e|m/ β���A�o]� ��uʄ+���8��'�B�dS>|�i2KC^�Eq��� �
G�^���O_y���޷{�f��ŹE�e�o]g�����FR����|�������T��y}B\�bK���B$�_�?ط �U�އ�SX���~���&�<Ʒ{�m�(oL��B?�].N�6v�4&=%�-�TV�P��;�);�m�9ybR���`X�"�	T����Iz%�NY�!|o��3��Z�j �����B|��;����ePW�J�(:G�O���2H���(aRR�{M]�3#�KG�%TP��6UƎx 愶]�M���	ɗIy�e��e���P���1�N[��U���8/�T�����M)��OM'"���ޯy fu�ӕ���v��A�w��?����e�+�C