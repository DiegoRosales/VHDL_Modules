XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�����+�z��0���助K>�{[#e;�7�uG����tZc�,��a>��mȱ+=mf�(���9�RM�i� )�F"9�� ��TC��Sd�y�7�Pl
�����1��wYs)Qe�3P]AUҠ�f��z�u����h� ����$�|����Pu��6���#��*���]�1n�� ��NPysx���lf����Q/댔Ι�.������($���)�M����w��`tg�{9Og�Ptҕ#4J��w8����[��D�D�ث��p��`��JP���\�-�����J�� a�4����T�^�K�n�?�	��8�ݸNz��t�A������&`�:K`&C�]ɺOU{��$���Z�m9
�3�G%�814H��+\`�0�ҁ�*�8��&���2w��yG����~����˵j;V��c R�r��{?���@�����`�O�,�cߡ����HQ�!5(�``N�fO��>���)o�k��{����w#W�V~�f������^�HVH��� �rI�����x��ӑ�d��N3%���"�9MMR�s!�K=;�U�F��	#6��ݟ-�a,k�Ɉ^++�����}.f����9rŊ�j�y�\8d�_(��
a�b���{�"Qe8F��#�o��0TO�����vrw���F�W�J���>��O����z�j�'���Vt�����.�����`cA/LqwE���6��ro?sD�9��Th�E�_��XlxVHYEB    4885    1380�Ñ]��м�<�Jp��T	�R�qY߰}�+*u���d' �-�r`l�0��r[�3gmjR�Kz\�@���f�h��BԊ����l�`����
��F��Yي;�Wq@�~��5a,$���l�>���nq?>�}\����]"R�AV����J�U�k�P��a�=��Ȗ(��*�>�Z�`��5Oj��9�FFx͏E��P�L���Io���6/�^�ґn ��|܉�l��v��3��
��mH���壆��)"��
zYn���}-F�� �����`S�o�WrA,as��V�2�R�n�q	j`>������]-�B$dB_�Q��t�_��I�,ݝ�*J�4�9�̖���>�	�cClI�+��7�O��Y#��}�N�#����"zv>GfՐ
���l\חv�ط�$N�J].�����e-��c�AX���*ʑ��C�-�7�S�
8�.�/�Ɂ�`"חA`-ѽs��'&�A~C�E�dH.�!�ԕI��E@:������$���?qN���-B�r؜$�XN$���q���&ҷ`�����b�J@5kV�^����n$[���2�ɨ{�zj��-��t�M/�v<�\����=n$��^����K~>��WT&��w80�	b�.G�����u��'6���&���&�$=v�>�?K-u+�WT��Q��<�/�� )�KLX�F cջ1(nPŒ�Z^ѱ�P�<�C��EP31q�fC	!6�0�
�ت��qqr�
�/f5��^��k7s5�O��q1^��Bݝ#s�i;�N���K��3�a�sN0��; �D�am� �~osڙ��;*9�K�U�B2���efy����w��� 3��^�������Н@
x��)�tb���3�-nQ���o�
?�v��0�ˏ��Q�<U?��&Χ���̙#N:�z�r��NO(g�>Q;g��Vsۡ�/��)��c�FZ�W>�j6�����
�]��Ӈ��<ڕꜾX��cvA�x�jl}_
�W�-�!T�o���[��u'>�>�w��@�a��P�����s�^������MH�?oǒ/\3�;9�-����1s�V�TJg8|+����ʚ��zg0�����сhk9�wɦH���\���,����qXXk�_��HǢ-�yA�36�!b�i�_��޽���ZC���^�4�,!�	��wD��e�he5V��C�����efk����k�\%���R�&����#Y��l�p��EV����_SR��2H�U���i�t7_��ӥL��3%��d��e�E;��$�~��3Z�������s8�(�	JP^�Ȗ����}��1��}�BS�����6�!�ǓA�Zåtc�$��cL�6_��~�4�Ry�Si����=�4�[pt*g��%����0SR�8� 4>�n]l �2}����4��x⸪�`d�dk�3y�ƈ�e�fW+�QK�d�\2������kX �O��F��?�h-�>[�����X�o�$ղ]^{����ۑT(d����?��Png�A<���m;����8	1�*�HT������-$�gi���� �.APWB}��5��Q��/ߣ���<�T�o��=`{��З�y�����F�d#���.���G�?q*2����!���u�����n6 h񠽫a=͛$I���@�w~�$L`E��3q��� ��z"ԕ�����!A������>C�sѹ�ws��Y�i�?��޻)}��&~�ߑ�Cpȋi%N�F(ӿ�8R��fYH��h�Fiz��de����z�[�ʑ�P���!?����v�X��ǘ&�c�>\$�(+����.L��Sl�%ZP�	\4�e��Q���5�}�A7���� u=����4�@��Z�Yy�dIh ������PeC$4MZ.�\���fk��1�K���������0���.& ����Kf�+ ��;aKtG�=���8�%�{�5j0Xgk
ǝ�"�w�����L툛���4Cgq�9���ʸa��/9q4"Y�~�ZaD���lg���S2-[�߀�C�0A�����+�G�` ��n�BI��1~!&1�(���ۤvL��;jmY.N�Ni[��G�5��C�<��r5J�� -[qG(6nl-@��c�@�C�d�}&���b�C���1gx��V{�\t*��-��`�S�)�})�C���+!�4ظSWX(i�6\XھX���ȋ{�z�~��,�D�����LF�k:����p��*9�T���Q!xJ���>\^�m�d���J�[a�se���z$�H��k
���ز�f�^=up7�d�EӨ����wyM>��ĵD���3U~1Ђ¤�����χ����1��fv{�e���h�T�e���}���f�?7��ʙ�5���1Ob����0��B�=���r�>`9k��QR$�*w�tt��}h!M�e <�0~s��5�V���5v�{�32�5��Ж�2�B��<4�o$�]'&�j�Jq�ܑD��r���-�r�Һ"�I��H��iF�K��s����wǣ4�R�Q@`bw���$,G��[S�b� ��{�t��F���0���d�!�d���Ɲ𐐃�&�Qk��2w,$�Ls9�
wA-�@D�#r�I�����f�E<1�@3��9^����H�t>������b�����z�,i0��3�Xy�\~|B� �N�{�æ��w�{Z��)�r��0m��惆S�����4+�����`�ڦ�3�K9�Q������u}.��l�aJչ-W��b`]э���.�*�J&/��L��n��C\*l
�x7ɇ��[rm���*.�B�ͷ$8��ⱺ�@Q�Å7L9,�Y	�
?�#�2��j�3�9���w�
&�d�ny߮,�㵺�n��Ҽ�%Ɇ�	)n�	j��EH	�/��!�V�߰xͭk�2�`�6����i���������^zˌΝ��RiI��M);S&���̾�Z�7�(g�h�evm���]G�Q�l~�\|[ځ{���ru7��"(HK�"=Osi���������������N��"���o&�|B��6��s�}4�a	d!9�Uw�
.VB���(�Nv�����FB����X|%͛���=M����7T�q��41z�ؽM��R۝O�[��}[��O�h�Z�8�5�'��s��!���9�j1�T���B��X^H\����t�n���G���P>}�5 4��a�܂*���	�?�C!2�RQ7���}�_�՚Hn+*�I:��pr2�C֟hPu=֕^v���nN��Ψ�$����]"V����7�04!H?�<�����S���VLuxWP��E�9H��"%JAB�*�Sp�N��d�E�x�_�_i	6uk!Sgx�C+c	1�/���m%�����"�*ac��c�)�]�\���Y���TI��&(�A���R��>vB��*���F ��G��V��[)L�㾋��k�G� �A��-�̯qˑ��-��]���B��w{����{���lh�w5f���p���D8�m�F4^�,��*%^�h�»/1�"��QYOݰ����A�k��!�A����H7��XZא5 h�L7]��G���d��ô�v��V��\��4I�ﯜ�)w.���J��~%��+mCw�$/���߂6Qt	��4���c���hW�ѽ��s���mE�.���s��*0�5�b�75Y�XG"UhJH�֭�,���pTb�v��J1[�"K����3�(�N�Ha�/��������lHZT��.��i��N:���Ԧ���򭱼�qwm'�kMڂ1�) <q��ڪ��Pz��^;��T��!p!v�b"�E�7Hz��
����)Pai4a���l���9�ԓ) -	=�f��J7�C�0Ե-��}�<sGyH��/��Y�>���>?A��`��H|�=&��Ǵ^��[ЄN���Vİ��૥�j~��n���w������#wg��ߜxH�� ��n�-(�REj�exxӭI5:��氩ҜPj(c�����Y���1q�p�?#����)$3�(��P���<N���H�� gIb=;E�q�Ã���a��O�H�S3�Q L�����G���.��PO� + ����6���~WbT�@i|>�r�ݜ;΋ײ��uqq�~\�5k����ܾ�8��C��1��EƔ%��|c��f�<�M&,]k��>�2��n]����]	��V~��bxTJ�}W�N�{	35�r���ְ�rB����� (�X���5I��9��P��AM�g~Oh��A��`�5�G{ �R6p�7��G%�Ę��J�vWfm��	G��	�j0qs@g?�?#�A�H�ꫣϣ���� �rY����ʱ���8�l؊shL8g��O:�0-r��r��+3��{��m���6���4�^<M�^�N��Ć���L��܇��iD��� s��OBX����P��/�2�.���s6�.�!<�X���o�s��z��u����	l�e2l��e����48��j���������a���[bA&�?�
�_?WR�S|�E��G�¢��s��m;e� \���`9[����]��H�]� (6d<+��{Rk�f�R'� /�8��D�_[����{���s$
Mh�]�Q~�x�u���879[�7��H9�|���J��3�w������4�	���2c�> �uF����Ͼ��ݻv��[��0an�'ÎR�8�3kg�!ٚu;�s���ެ7�D-�e�����G!5|S"B�ZU����O�2�4;�/�r�tW?�(
}�W�s���n��G*Z����D����:���q6��*������r���IIVfk:F�up!��ʠS$�����*��ٗ��)�,������[�糰������