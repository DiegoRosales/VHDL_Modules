XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��R��`/�k��W<e����m�1��wA�ǈ��f�����+,�<�`]�?�ZEV����TWy����j"��^��|e2Uu��ȕ)��������2�(`�.v(Mi���N�"M��D�v����~l���W��y\$�e����Q�;VJ��h�A6e��o�^���,���Tz��������C]S�#:Zm_�;���޳X��|]�2u4{��U��T�KI��w�:��W^�(K�����(�U*+g$�$N3	�m�OuX�0_��!`�Z [���?>och)"H�'���}JKT���ɭ����4o|�N;���v��ip��D){��P����Ϥ	��Յ+�;�ݼq����[�A�݉�(&�& ��<NN�(��U�����eʓ;}��h��%�E�L��OkI�|!)P=zvwC������v���������� �8��~��)`��8�(� �h�" �b����}K��v#����1a��.�wq��r�w���/�Ֆ��%��sH�U����(@���y�SЯ$zLz"����2"���Ȗ��[��G��q�r4l]d����q�Z�����ƅ��g�#	az2����]�Z��;�Ac��C5���B�g��4�ⅮʒW�uB�FG!&�E����WС��~�1��̧v�
u[�ǣ��y��� �{��ntL�6�B�����lZ�j����W�+����SZv�)�&���bǶ�=5��&-f@Ӫ�!�.�m�W��X�M?�Y��O��XlxVHYEB    80cb    1be04���� ��U�z l녷`[r���ݾh;�KcpL�ܛ��͸�6���9�~>�
����J7�x2q����b�����$���ջ��LY���yN>�y�p����+��Qԭl쉅��e�%�Q����_砤�{i����9�Zl�U��I��Y�����z�?�ȕ�8����X`��΅��1\�_��bQP����iW���Aax�*ߊ�I�i�f�y��c���3B��:W�N�f������l�kp�;�)6V��u�'nkM����pM��a;
�WOX-�����7�7G7iw��!�A�Δ�ذ� :8�s�鹡J�vj>h��}Yj�.G^�׫gg���ߴL_��	��Pq�UK��$���o���m}2�g�*x?3J,�idj��#��0��*�Vd
�*�(7�}��r�C��$����&��/���
�%mS�v#2Q��	=��Q"� ��F"�dQ�7q�qi����F�A>G8
5��R��X�����Pu���[�9*�
�Iز�^6'F���­8���-��!��l��-���u��X�v�җ�-��V cW�2����wO���9ea���~��qu�_?���O���X�_��!�|P����}�`�7����KDb����Jq|�Z�dyQ���6���omoKg�cc�%�QJ�ǥ�Q�siʟ��w8���X�����c� g��/�=�=��5 9nsI���ƈ%^��k�����4�1��05��o��e:��/?����<��=���rQ�3������<\l�{�X!��!n��%��͡R.�Q�$�j/5N��1(��������0����*���P�]c��u#�<��1�� ~��I�X�$��ੂ�	�����<4s���c�P���g�6t�k���F*F��'P�M����@��W����1<�)Y��7����9�DO6���i�P*�}��/��m��\������ףʅl�
sMGF�MR���ݐ"�1?�������[�A� lE�j��nq9�| =ղ~�ZV�g �s`�:3�P�Y���K=�KGo�d5�|��W:���7ՙ���h5;�I*#X_� �Ib�� ���W1�M��5
j�h]����ȪZ|�G,O�O����I��g�t	�5��lQ��eFފw������E!J�߅e��vlʣr�$��U����K�i��"�t���#6�ESF�7��	
F/V� B�v#ho�|2"1���ZS���3���~*�_ �E��ޤ���C'5��OT����א���5�UjVk���I�2�>iN3��#X1�.=�ő�
���FI�����n�"�L����Nn��$�h[�0U�Y�H�'h���1|GE�����׳��Plcѵ�G�����T-�p5���Uˁ���b�'��7qQӳ�W�KO�Ы7[����ؑF.K�)�UI�5)�@�_6�z���H�(e�,L#��� ��n�> ���po%1�ZB|�9Ǥ�kQˡ ?&�#��z���hz�O���ͱF��-��q�dl�����ŢM(���DS�������mz�2b�kN��>ju׳�#^�5�a�$|���.UZ���4JVe��/�
�ܓ��/<�u* ��i��/�m6,y�;��J��B��Bb��;pJLY�p'��Lb���(��D��2��V�,�x�G��)���~q��{�k:��Rد�<�
���	Z�؇��1$�űt�^"�&��D�H�A�B��QG��}5�uf���y,�,�̉�&�I�{'�n��rë-	wҰ� ��L��Z���e�튣�NV�@����I�d�4���`2�E������ �I����>�ӛtH��ׁ�W�WߡA��I��*����'�g�wQ��`^�f�LViɓE�0`P�{����n,83�`? ��E�?J�2m���6B��]W%N2��XA����v��ya�X�x8�J�N��p��!4'���V��4}263���a�� oU4���iHU��ȍ�F rx�;Ơ��jb���Z��&�nAܒV��Cn����Ql�}h2`���'K]�� �2U@���.�#�k�,�D��t�*�M�]��)a�ߙ�}ê6��X��t0�|�o�i����8���e������#�2�1�0JL���:�)$�K3��e��?�7��i�.Z������]����v4�U��6�_#������M�[8��.d�O+4,��ۿ8V�m1iK��p�J�|;��ZF)@d�{��.�^�9�7
��	���N�Q�=�#�Ԑi�[l"D�#��L�%��$P�l��b������������bO��A�">���s}=�,��-�v .�,dgZ�l2z&Й���Δ�H�L�p`{z��i.<>�O�_p0p�K��>�yȽ�3	5�+�C�
ե��93b���Tf[���aUi�_�G&�ݲ�QK�@W�K.@}b��;��3�w��P�
�� \ܭ��J�J�?	2��X\\z��}_値;u�/��gh��;�BP��-���P��l�����`Y�����h*���/9�n�N��^{X1�]A@`a�R�qaL���_�2ՀЊ계!��h�����hl��R�nF���ݘ��-=<�CDĴ�\�#�o�Q�W��>��� ���OY��u=��bēp���]媼�x��F;����rǏ��p�f5�����6���A���ckR}��f�d�(��f�7K���-JM527��&lo�[�PR7��J�U%�YK������������ i�������x��=����%M>*��iϾ��)��.�N��H��n���-�=q���:�jw!i�%��u��FN��dǽw! ?��n�9z�����b��j�Y�M���q� �?��+�#n��J�z~.�h��t����.�6�xIW0Dr�.��\AD4��az��͈>�ŕ`���*�X�Ñ
���J�,��U'�G8�N��+-S�+��X
�5|o�Q�����(���)��.	������E%��i������f�$,�a���1W�Hz�s|ϣ˯
�f��4�YS(��;_,?m]޽�F���1�|S�va�҇���:I��[R��iD�'�C��O�~6�@@�����[Oԃ�6d^�W��xb!��c�������t?��䘘�7`?Dh�����]��D��F�{��P�o0B�&�s�S��f$�| �^��p�r۽_w����L�����%���0�7��A$�r���bn� ��\*�D�Mceg$�@Fڼdu�!�B���6x�����+��f�K��̝`��G��f;a�"l_��ND.���hw�������"O�<��h�z��Ѽ*T�N�^]�0��"�[ϖٍ;�d�w_X�6A�F���ȹnM3����G�-�9�����N�t����@:V��6n��.��)��=:=|���rJ�9;��U���d.�:��]���"�3��T3�h�T�@�1�W�\��yP �n�}Q�zM-<}-#�H���ٹ�r��y�s�c�c������`���U�K�;9��e��;e`XHR0*߼�R/�5Qj%8 �{T�~� (�O�3}M���l]$�ճa�ǝ���̐G��%	���sߡ~����͉��0�tu.}f"7��r�=��ZA8ݤ�k�&P�wE;��xo��G<��5�hUo���}�Q*n���6���!�ίu������\���ݫ����/�r�a��F��%c�j�{��Q��c._�fn�l"�er��r�V��/cv}�!vPl�O���,͇�j"��)J�GG����7,01�*!�W���8� 'L��h�+���"��c��R�t��ҔP�?�/5rU�u�3.N�o(�cҫ�V������H��Ү�2jGrq��~&� ���ղ^������i��jO�oz�J^,y�x/C,z�D���P7�"�t�7�֊RE�k���.2u�N��ѿ���w	�1�{��Ėդ�F�Z�?�)�}����,��ҤǢx4i���L2��"�� �kh�������5�)�˩_���R����A�A+�(q(!��s���o3τ�j���@�h�$a6�9/��TbnE��AS������^z/��xQ���~#�Q��Q���n��t�r�.{���*�t�����d�^gU�xR��(/�Fy���u�o��s(�B�b?�� 2��+Z1�5uM����	��Y�W�~l����ePSE>~�)&��nA�Sbb�����S����UJ	�ψ��^I�y"�W��7����j���䤻�e�]H��-�h���b�9�{������cf���
�GA�sj�Z|�% �B,2�U���WkE��\1(����a���f3!�kN
�Ȣ,Z����*ŸO4<�ġ�ڛ�a����M$�Ǽ�������ֿ{W�n���Q?X�"��'XH�L����^�%��p�qvA�̙rW^���*�z]'Q�N��e��=��#��\�9��C�u`���HH��l��]?L4?���M@�"�WO�1Ō�q�GU�p!��,�)�1H�����Z��s��v-E#����-͓�+m?��ҏ��/D��X��=m�ق��T�\s(=�
�h\E�N{B_�C#��hk���(Ò-"�2�iG��*%���u�#+�D�-�t���O��E�g?SKw�s�D��~����0�H!4�I�}0���~O��:��s������dpL���O�a�
��������@�PM������S�St�9��&^�
_���5�� ZY�G��ԕ7��H	����/G'�`df��-�Е0 ��G'��M�4���F��}6�*G�<K����t�/A�U�,B�ķ�����$ϯ2a�g�(�/1f�6bf|�z�A�ۘ�[��eg�m�����oȨ��_	���4��M;H�^��t�/���.�6�:j��}�����|�Rf=l�*�g�˶��=d�op�%��Rr*�f�����]�V,����S�hLS8�TUa�kdV�<���Ґ�q8�q�L��^U�<�x�_K@�*%�пd����5[�� �1`�`N*7�|pڂ@���un�A=�0�����������l��P� �������%�fQ�b�_��\WZ��H�nO�b�&�u_�^r����˛�����vy�������j�덀��O�W �d��
��Ϫ�����}P,'5��s�{��F���#(���kY�cW�u��n��Y��&��J!~���m���VǮ�ҽ2���9�5c�XH�o��'��`�[z
P�N�jg���8?��� 2�10�I�S�'ec�ˊ���.>��E��G�`V㗀Rǿ��j�3N�����q��{����)��z��À"n��Oot@��FNŢ玙n��`j4��r���@�)RC����k��\z����������!V�{�m�m��θ��p�*3�tCl-EH?�nw"qKH,�?Rl�%K�i&�4�o�K�+��ނ�}�nD�P��S?��*�7�$�S0����D��\�Dd�-�w2��T����ߖ�"��cTtݜI!Ⱥj
�E�н����͆Y�5�d�!�|�lXf����l��.����EfMCC�[
A��팥���M\R���T��f��nS%⃢�OA���$���]58f���,!}�}z%�Yx���-$n�i�n�Ob���R�!��t�(_�'>�'qnd+��w�Cm���hu���.��v<��]�f�$"M/H���R��$�>n��H,cDLO�/�2H>'�|~'���b�p��߀�#�=��v���%p��m"#	g&����Ѭ���є1�G7ƾ�6�O�EC�JI�#�L�(9[�B7����|u����z�?ع���gM�PԙQ
~�|�3,�zo�D`b�`[S��n�J�b���	�Y�L�\�;������je0!�%�`܉�ȶNk�>����:��B��O�*L=��`�+|y��薝�u~`�EE���Q8!/IjxZ����Z��I۩��)MKM�Y=���ȨWUr��"� G�Y^�1�U��-�K�1��Z����7[@��j����!� �ٮ�r�])���]�� -�}E��)�F�_�w�_8w�-��+�#Lh4��N��|�A7\�y��*%y���D��dy���V���d���kC ��aT�3eˊ�� ��1�2��9eo�����颎�j��7$��G'�:o�]��%h�'��UH��>e���%��������{��'��a%������Q�-p�S�̽:ܔ��R�%�\9�%��^�Wm�Z$��7(W�7^Gŝ��_�>e�gb��"!��9Z��m̫���*��	��X3�>�ۊ�~W�GO���g���rt�>�d>s&nSF��t�o��Ν><�0F�fY��(�g�S�)��_�V�	��jĂ�!.5�L7��RI3;)Ј 	���l?=^!D�L���|����#_�y:��:?����Xs�Ms���Ev��!���A�6����V�/r[��X�S>AS�tjd#�g��Z����T֣��Em�ϓ��Z�F�G�9��o�Of
 lqIYȫ����#��:�H]��Q�H�5�I*��2�`�d���v;�:�EMj��d���{��B����Qآ�D��g�0�����:U����	�L�_��I'!�)��n�@k� ^��+�7�z�	�oS���yn�$,|�9��&n �O��G �����y\��������j�.݆�7:Bm��*U�5���A��5=.	��t	>�A����5�KFRr�����p�Un|�x`���+�u�Q`�p������6p~s���/���d����.����B�<�Q���yJ��j���O�`xn�4�Kϳ��A���A�aY@�r��e����օM蟥�v�h���r��=��ӏ�U�dA"2��������`��t_�A\�H+DxU�ڳ��