XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��+����*U�Y`M �����:dݍ��6��=��%�m�Y��5:+Z(�b
�]�[^����Y�#�\p����U��1]�zc�UF�QA.���ؐ�����Z�����ٶ���_(Y����Y{2P�KW�B�s)G�]�����{�)��ĸ�H!#�%�Hf�p����:�X_ 2�U� ��1Ē;�<��Ve)���eRW��p靚�Q� pQMl��kbP��e�)"[���^?��n��ٻ6�k!�K�1�����g3
�	��z,��1c�ğэ�ۉu*\�1�J���eE��H/��S�ɀ6�d��	�w-I�ڕefߎ��Vg)Df�
x9j�.:�yɢ�2���'_�5ԓ���L,�P)Q;�ä'%1$^A^YW݀�\PAG���
��U2Ƥ����N�c�)���Sl��o������6��$�zZֱ[�5D�m���y=`#�qѫP������ ����x)Ee�߇Ū7����8#]*�FB����Zd�e�^�c3�3����s?I�,���.��gin(�w�Jd��Z��\��l�u����g��9k@Z�zB�M+ȓA��k���1�\;?,&(��ޞ��I2��8��S%� ��L� N��=���Ç:H�.�B����hH�ƇYE��amBMYcX'�H�ģ�Ga��K��d��sF�n��]T)�]~�<f0����
�ߐ���4�`d�N�W�s�����.��'�H��!�Ns_3�CT&�<���%�{XlxVHYEB    2962     bf0e��\|:Z7�dU=r`��i��_��;I��9�v����E��7"�ו�D�е捷��6��Y�D�!���#��O��S�'���m��߇;�)��UqP �ffg��;=dP!R��rM4K��`D��!��8��BI	U��%��%DGZ�$��)W�4��]�܏E�L6��p'��#��qB�̀�� I��z��	,��t~I�g���C�s|�$9�U�1���v�i���z�M}���F�G�r�"v!�;�?�������1�#��\i�o�4
�kJ���J����?���K�;r6?�3����M-ћ1��Kh�)�զ�|��A�vD�HG� /�T���|��]�W���7j\��N��,�@`���#���]\�J���Mh��6��.7*�:��;ޗ�RJf)CJ�xP��^�b�ȁ����������tc�=��p�:�*�����K�j��[��4���=2�N���Y?�c �����^�=���AU9}�����ET�!�6�F}�r=�tg��V7��{��X'��az�/�JFβ�Y��_c5�|���mi>5_?<�Л�,�tx��ei�ّQ���y�Lm)T�tа��=RE����Rs���v�o^��R�v7�=�N�tȢ�����2@쁴��ڌJ�����'��rH����q`c�W�>�x)��EY���:Sx�2#9��԰wp�%jP9=GgJ��]�1�2��Pf��J
��܅�	��땔�� �`!���6.�𷵻^r���7A�����š|A%�E4�/����Whg �$дȌ�#�-Z�����(�'��ggK��]���-��3������G~���0)��0��3X]��Vӧy��`��X����|]�$bNX�l꘢�	�s�����6�I䅍"6����>���SP��}^LRKO��x<��d'��]�(��.Go�Ԣ��;vi��sq��%��{2�c ����`�q�Y�`�n≂�߿/;}�"��h ?Q�D��j�~W��%A3���<��g�^�����R�*�U�ͳЀ�G 2�M�%��U�O���@�`ߩ��d9 
>��v�Eh��S����a�lvˁ}��e�u@k��{��M<����_92k���EL,A����,(�"�H!9�=�+4�� �w�6c"�)���춧�2$��N�s�t���R��K<����� *���xi�ϣl����`WC��R��X��e���Lr�!@8�Fi�#�Fԑ��ʙ�����k�M��3=��ſ������9�52�K0R��O�3��9!���G�wPP��*��<�6�8;�b����4HP'��g1&^U��j�h�����.�6s����R�4���+��	TS�P���$��6�P|9O�Ty�Ic�ii��Y�1���Kս�~���3� ���eY5sQ�A�,��"��3�q��Z��齳����3JS���+<�s��`3qW��j��R�s����7{糸q�e7�Y�d�Ӵ�ry�m�����5��4H|�S��}�����q��jA��'��lFӆ:��C�D0���HSM�e��nM��TG,�A�!*8eA���\�ɴ��(C>��Pqs�r�IA�@#�G��G>�.�8n2+�]��=��1��w�B������.�9��@`{%�}[ca����0>F���res��Q�/E���H���C�d�(�4x�i8��Өt�e�4�NM�M_��Jٗ7Y��;Q���)4�/��|z�7d9ܬ
`������-x�t���u���k}��*]�e���Yr?���p� T����<4/�`��r���[r
uZ����iz��g���<�q-� R����Wͯ�[�5Y#ԡ�)��(i�Dqo���'���O�0u��l�>)�^7��]��N�,*U��#0���z�H:�Lʇ�{':8�Lw�K�e�ߧ)[�܈���֮��T#'�����Ԍ��bFDcV[�P�����P����^����ȋ�@�XP��X������lGj��~- ��ڋ�x�BC�f|�9\��u&L7b;��k�0"p-�^Ճ�S���:67Xn_
����bc�`Q�������\��T`&�&��%&m��h���m��x7��x�F� ��{�]x�!�LQ-�E+nSn���o��Nvٟ澗��"G�|�������x(�G�13�/*l7�J�P�y�'y�Lb�k6ܞ!�A�}0���O���]��gm>ǜ�w�������W��f��-���~W/��,l�ά�^?�(��.[��"p�C�aۧ����F?��i�S�G��T�Lf�=��eX5A.��t�-2	..0�$b��Z;�}��b�j�T��*����"�]�Ɯ~��E�%���M�����(ֳ���th���2X�ҫ^v;:��[�U'���*m��,om~���~V]J���
�O����E纡�m,�GH���u�aS`�ӏtW
]�,�rUQD�sv��3Ħ�T�f���cy�"�:p9$���"�.��ݪo���e�L�����-�M��y�C	���e#�/%=��2�!tз��}��0G.�vx��ث�O��GyA��޳�h� G�UQ�^�ՑQ��}�V�?&�O��S�����Z������������ld��]M���vX�|I(��[��̀&�3N>D��15�8;s�`�հ��P6���/��	 S�����~�8��DK3��k0k-��X�q�fvW]�n	a��,g�F�z��oG"f�u
��j�8w��^�4?�a�JW��*K��9��R���q���9�����fhx�-4��E��6�# ZӸ5��3'�� by�D�{�������GC���s� (	�w$��^��������]��ٌ�C�Gt]��ŻX*������5�3VԳ]5Ѩ�_���*l�6���OO1s
t�` �`����������&����F}i/Zw���8h