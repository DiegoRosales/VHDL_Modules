XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��.[h��z:�*�䐭�m{��޲|�o�N�YwO�+��}T�|t0+l� k/2h-Қ(�$��4ث��a]�pw��{���Jf#�󐾃 ��#�,�Y:�`��y����#u��2ǆt����3�U=��;�G�|�03��y\  8яn�p�	���aj�ը��d��[��`(�e{��+����	�J�d��W-Ĉ�Eq�8(�|�ػп#LGqN���D+f�]a�����T� ޴���L@��"}x���v���3�M��e����sf�h���0�Ms����yX�N-��B##��w'!¡�Ի��8C�'�>V�!�.2;��C<��OBD�M�����R��50_�^k �iG� �^9[��XKc�q�E���/=����ʯ����?���s�y"p�0�L�G�KjXU �gҔ�V`&u�Z�%|CoM6�W�u��Mt��ľ���I��։���&����R�5�P�ӭE�^���n�r~l;�*Wx�Ծp�}��Ɍ	����&G]�H���g�R���JB>�6t�0��*L��0C���l��`k�w�[��,d5�*��5�N�I��0,ɽ�9W�rP^''Q>���`V��iG$,�����-*�?,h�c
���S[�)N��O�q�aX���3� y����a�5���8
pК�AA�T�M�>��1G��X��I��*�`[D��d7�׭�9䦮u����?��`�!�����Y C���A��-Ԙg�֑D̟XlxVHYEB    49af     c70��!�N�tӴ�aP؃���1�2�M���Nڄ����|�B�G����m���o�](�5�^\���(�W(n�ѵ�<K����� ��B_���B��s��f�O߼8#�S������ޱ��j&�x�b��٣�Yy!��WV7r���9S]���iW4:��"Z����~�h\�=�|ݓϩ[�Or��uV�_����ۡNQMi�ߤ!�����^h�"Q&���Ban`�5���������w�*x��A��Amu�T��{ۆ�tF|,s��ś\6�"?a��֗��K���+�;�ѷ����j���));x�{eC�%��k+1̀��
�����Nه��/	ޕ��'�j��n�yf�r�CUCd�'�g����qP�B޹�כ�@U\�����t�D�ا�M�؜�k�UoWi�S��O>�}����B�$'s�}�y"񷥰��㏏(�h�v���3���:S����E����iֵ,��US�b���67��q�n�>��y���F�Q��6x��PQ%b�h�ꁖ],���*:Cj�oO���5�)�\�/��<:�Œ�t��1�Kx)Q	5���WEǾfn�8�#�!�FU~y.l~Qw��C`�g
S/��&3A�3�ȰX��|3�� 7�DăJF���U�UJ̺NVo�����J�x0�p�}ybf1WQN"]��|�Z�f�K�6c�8�^L����:�g��E�J����3�<=��v��y����$��®L/9sXV��}�*,X�q�Q~H�N����f�u$���-(:�K�����J����H�r��͈�Im����z�^��!jꌦ,���|�}�#n�:������~�+�P�{����[u��c�M��Ͷ��P�[��wz ���f)ZN��E� 暼fk��
�����6V�C�� ^�@ى�u 7�d�X���a	������T���n>���#��~�ѫݵ��9���V����zH�k�$Z~U�Ye�6����o{���tp�Ő�=I�l���e���rH�ǵ��Lǻ���u7��e-�>�
YR#�?�k�!h�w>5d�]a���rN^���0H�yn��$YSvh�c�9�/�?��'��l�r�Y�0���?�YH2��W����eӮ� ��OU'����qH�nu#D�h:ߩ��C�'xߞΖ�ְ�#z�����\�>��ei���m4F���8JLο3�]�t�^��N>�:��]�������>�^r/��Ol�N]ܞ�͐��Ru��aF�p_��-;�ݶ=P������l#M�����I��i������j7O
'o��W�$M�#����'��I�Q�m����a�ޚ�5l/�{�����ۡ0*T��ې�՞M�A��xk����7�b�X���������θLPPl��[��NW�B��U��/���7K��C����3��Q��ii{W"����F�+Z1`oxD��Y��<fp�Z�ϋ�<�s�+1
!�w�ʷq�����+3���u餔 S���?>9g�����ޒ�Q?��n�BJ�n��y5*b���O��dl�	��
��&��ĩ������qܦ�g:nx,�]�CC�s���ö�N�'�̀��!M�v@��/uO.>� 3����hV��D���	��띆��<=Ƨ��k#�����P��i��8��ٖℙ'*��T�6�Ǧ��	�B�����������SQ��KPz�uU7��v�	1(����2����Zו��9�����5�%6`����LPؽmU��:O�wW	�>�4^}����y�������\S� ��7VX���Zq<@m
U~�FĻq斝r�5�F�P������7h����� Ѫ�X����j��M5�F��N���^N�~�0��+���k֥���Smfµ���u�;5��K�G�S� �� �X!�D�UjT����3�a�k*��4�܍2{�����a ��qe[I��4���0�AOی�xŖ����>��*Ҭ��u�
Ol���w�.X�y"N�jn�����=�bap ���3>Y�l���"�4��x]*�=��� }����L���>nT�-���.x~ɵUF��s����u2LQ���yxݦZTt�-�1ѱ��fsU"��0��b_%n�E�D�@��VaUJd�f$�k�uH=�k>K^J�B��c, �]]�ܻ��|����Г�t?&�o;����އ/X�m��
�$��WA���*K<��`���
����<]���P��h�A��F�B,��蟴Ѕ� /S�sps��.j��%����X���{�E�
^]�L+�*\���@�*k�� �ʿ`�>�Gn�[����w��Hv�2��%���Q��4R+zRۥE$ v�<h����'E��pk�O >��sBf%ͧ��a#8؂s�'Ǎ�ukJ[gҥ]6����/
�)������|v*��Ӭ�?�N!/�AX�����eA����'.�{�K��U�;��.�;�fT�L{�`Ы��8쌞φj�3��r��a�6��|\S����T�W���N@^�1q��� �z���y۹����/"�7g�k��^�?�_k�W��_J�t�qt���Q�)O;>���z��'�j�<w��`D'ΠzX=\T�\E��b�ߨ�v&�͆�x�+�-��ȝ�uIҢ>Wm�D�'�:��{�@����C��v��ȩ������*����	��'9�r���4�ۃ��y�ď�ɒ)[�>F������]�~s]^/�ۏ�J�k�^lj�j��N7��Q�?*bb�oq���w!
5�����{b�j�b����H�t����0�Q��Ң��G�Z���y�3���E��c��T���;��;�\1��;5��0�S\G����]�fs���6�2���������/����^�/&��Eˤ�_�9���%��_�z��9]�����v��|��'�E�n�ܾl���q�-a ���E��JMt�@����_�5���5�οH��~�k��&8�d����ϊOP*@6ȡ;��?��>�=�FIuAs/39��+�mMr�=�����F]8�1�);ƜVa�h�ӎ��G�C����r�ȅ���w8=����=yЦ�S3q���7y6