XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���S�5�\YWs0�9����
�h�Z���;'+��{H�s#_�3)�z�Ql���}o���X� �G���'���\Q9oj�w�κ��/8�f�t\�q���-��j�sw!�Z��i ��D�alNPY�r,�����ޣU.�Ƈ��t	�����T��IeT�A<�m3Ζ2��uD
�a��m��h�j�eQT�yu�M�8��k�b4d�H Nĥ�천
�IG�Rk��-`"g��`{|��	أ�+�Ɂ4nƔ��!��u�{�a�ۮB�������yxX?LԿ���MxK����\�<߯Ҝ~_I��(�ʧP2���\�px�<�Eϳ��ĳ/U9Pd+�ۑ �Q����Y�W�k7W�Ԍ\6�(�y��/+���6�)��È�=�[�&�8
Ʉ-���/�iL��S֡Z]�w��cw��?����8B�w퓙�C~�P�c
����@2Uﮉgy�ٽgt��GDH�:�üJ+�(jq��[�2H]Q{����(���8J��M��@��J����Q�{ư�P:��'�q�����2�(��T�B��u� �	m���%���f�v�E�8�G|%I�B59R�1�����#���~���y��ة1�R��T	�������� �J:F/$����αh�k�e��9s�8�-;��ѭ��K?|�ۖݍ��H����R�h Q�㺕>��<0p���Wj���n�J+J��7�E��O@=�_0B�!/��޸�}�q���53��XlxVHYEB    22f5     a609#A(�����ɟX�����ct�hFUx���}�eP�>���2��Q����y��h�5&���ݳ^x�&���>GpɬKp�g���>Ō��������#��=����]��L�l�a��,�a��[p-q�ER��S�%������C�����O�'#V�Bem�h��\'���)��lC�����:���v Ӿ�#D%
��D��k���gC�w���/��UEI���m4��A�!�����ӭeX�@�"ā�FN%�x�h�s�,F�0'��n��n���Uc�<x�U8x�ܞ�b��������?h/ى�h�I�L���0d��D�x��
�"�bzI��مˎwBe�=.���V1m�M��K����_�c�	9I��P�� ;HN_�o\߄O@R�`'�娹� ϲ�9ft�N�������i�h��&=�k�''E�+<\���Zd"H�}����)�$�<��c|�e�a�<�k�0���:��7��3b�N�����(�������NR������:@�������h�C�ײC��#4�6pɘ�Q����3@��b@'(�/�Ոc��UʝS�f�y�;ؓr�
���	�/�kP�Q)'��Zv���
:\������ѽqC�4�5��DN�����!J��<�������U�liƪ&��7+���@���g�N�qb$(�� E���y�������^J�� <Yn�9m��gHZ�^~^�
�뗣��>
��%-�u~v*=_^N+�Eu��0�����Ь,�0?Iv0�^�
^0�P&�\�"��3����B��c����`G0�J��$�gr�E��>���0�^(��x(�/Zo±C�o�@�V��ƪY�5{%4 U8i��T�B%"����h���wĤ�,!��{�ݓ��BV�A�-U�����_�h�ϝ��0hb�� �4"��Ls�03��-2
d����r�!�V��SA�9d���b� !y-�Hú���;t7����h�\��=� *)X�`������W��Q,�d$ؔ)Դw��]�����s��؎� �(S2;��>�~57��ӽ�3���0�M�B]+�ЈiK���������9�[*J>��G��vp�i������´���楇i�ޙ�?\����߫
�$�������LS+�"IFLj���נA܅A�.�듂�,z�.��%�xB%�R��[�&�����O�L��m��k��y��W2�sA��ك {N�GnC�y�4���Ӱa��G�>�Z+�bG�5Πۀ��و�SR���Lv�>C!�]�lR�2x�?�2���2�|�^��y���Fv�W�(��N�� nY�ЬB`x��N&pn��1�\sDQڠ�x+�s�`F�C�D�&�p�xf��'L������r���)OW�c#��>�.s��,�B�6�RM$z�*Ⱥy��A(E�P�G����*}b��Є�f�]�����6#*���3��s��0��P6(���*5��<�sV'�0��<�4:��ImWiϧ%�f'��2>��}Y�C�jD3	�ީ:�P�N�$�	O�2-���vv�����pn��b�=��AXcȰ����B�H$��زqZ<�L/���Md6���^e�i�~�7fډ-\0��i����h��}@�ڽ�仌�y�v ��V�dg���(�s�9��6/y.�x�3�9��C)��T��Z�1�γ��T�=���N�C��e��,�x���|z�|f�R�$�R��>��/0�_F�O�p�d%�¯C��)n�4�qW1鄩�r(6?G=n�^WW��y�����m�H���`���g����ί�����L�+�`�������DS�Xҵ����j�V�qx������!�4̮|B��.�":7t��(zP����m������֪?�����~x��%��~��(��0Q���u����]'x��$��Iܳ�Q����:�{��h(��y��-B�-vE��;��B5��lUY������:a=�ֆ�a�n1���u�Fc�1�a�Y�)+���_�3��Tu��z-Y>1@�ܚ0W�#���XL%F������QB\_�3}�o�G���T����7�t��*�'H�"g���ctJ��<�y9��e�3d$a�Pj�I+0�b4w���f����
.��X�(�s��]�Ĺ�h�Dtg�*_���eE�����v��)\N/P��΀�i��6���8��@N��2��rA4d�X%ӈs��.f�1$sߌ5 ��Ybs��� �{�xaչ�6���ҕ�c=ν_�nC�w@Y.n�~^̟�Cx���.̮ϻ��C���hxb���!��Ň���'��姛?�� B\R	�������_;��E˸�ł��Sՙ��$,�v�Teߪ��j���Զ�LY��V�0֍��J�A8���]�I(���Hl�Jp�7�aѿ4��Lژa��>�eS&�m�P���V��"�(�4V1��߳7ꞯM�s,���	F�9��ْ,l&chZ��)}n��2q��E6���{8��5��u� /{>2�P����x?0�!��3