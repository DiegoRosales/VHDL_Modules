XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��}l)іNk������~>�Q�) !LΩ�(�/�g�t�ѱ�����I{ d8[`�ҫ%��x�q��*��B�Gn㾆�܋��3�d{�0�	�_/70��qW�z���"r��i.4�{���2�2S�qZ���i�7V־�hk��V�嚵��}�ӽ����	��X �-x���w��gwԊ����m(��kɲ@|�Z"*�Q�[�����|�[�S�R��l9g+�c#޸�,��>�����m�L�$�����8Z�����x��܀u��T,N�z�=�(�"!�	���SV2E{�
�S���� ��� @B�à�~"���ՙ?�h�bA4��%�|�s;݀�%i9ӳR �KJ�qmdY����E��[�;��X��<���Z��y�N��_72� �Q���UJH���u��Vp)>iڛ^d�0O����܍t5{W3��"D����D�Й��:�nD��n0J�hq����R�D���2���z�yg���[���L��1eo} ��<�nu-ϫ�mV���G�z�(���(�O��N
lY�.���n�1���g��2�}��Z5�O�\��ѩ���h�J�dh����E�h��d��MH��P����[ب)�\@P���$�r`#	���z�bhg�ib��6�f\Fv|4,6����ԃ�D���#t���nςb�E8�����M]��.�������+9�s���:F���dō!��&<E�
�U�VҿFژ>Y�?e!�u�l1'�nx�W�iVh��@?獱XlxVHYEB    30ea     ce0ɍ\��u�+�0���i�.��1��B�?:bh;����>T'�8DH�H>� ��՚�Xg(g���p㡀%$��RB<7�Ok�pkB��f\���6�����yryRٓ5,�τ_��=�:gp/�ߢ�ER`�'�O���p���gJ�H�w "'Q�B����7����5t�-���o�J$�L�.��Cz���\���L��F��P^��L1u6�E�.g/өdi�I[��5F\�}g#�Тv�Y!�����w;ܣ�٩S��=�_�(��?�^��#%Ft/��~ګcG����_��J��S 9yԸ�"b���ϰԮ�U�5m*��%��:w%]6�B4:/�l#BP9%n/�W�$�/ԵA'�[� �E��
�h��%�����'?��R��?fB"��G��|�Z�����i��c��{�%'=eо��vs ��HԦG��3�u����&�ye��6���NҘR�qx��!�I֨_\��ͭ��Zw��!Ic�\5E���h��gK����*�<'S8'��7���k1�~5�}�3<<����/((�B=�3(_��|b��<�����^��|��G�܄�O�9*�w��%�O߲>�7��k�����p��v�,e����wUWD�0�[���+݁�5%N��d�6�E�ױWq��r.^HƏO�8�a�0��ޏ���<#��H� �.V�H�83\����8�o��|Z0�J��};��^�Ju_��˞G�7|"���ʒ���t�͂�����~:|�yvg�Q��˸��Q��&������!�е�Ø�˚�F����ݨ�ϖ��L��C� �IwtB41Z�BS�L�=��n���u�����r�U��[�>����h\���y�V�랈^1�[_:���ӭ��*}���/���*����/�G%�g�pc�(!�4"�}��	��e�4"(�+���6Y<ѥ�=��ͩ��?���)o� �`��78R����h��ړL���ÿ�v�	�l�?Hd�5��fk�&�1��+$�v�R"��Kc���P,^��M:���$�GY�2�cJdfW5Iu`h=��_��"͊�E�E�ϰ2L���z$�=F��O�݉��%1�gm������z߄-� ��s���"�1���V4�> �>�5w��W�Ѩa��U�#�H�M.:$����zU��[B=�޿�!�.�%���l?͎��~� �Q��ҧ�SE�/B�.4�z�F�M�!�7"ٗq��7�^�5��r��v��Ij��.M]i��4�P���.|�Q��_�K+@�Q?M����ض:y��{���NJf���q�2����ǯ����h���e־�x;�����ij..H�[V�wU�H�?HT,3ɭs�CP�]1��?� -���ͭ*_M��F���^��ҦP�K���,dx�+rK�wH�*V�XhGV�˸!S�e�{�y�ث��0�3���MK���k�6q��L�#5�^?�<�d�H���Eg��s�4v�|�2F�}.JM/�5zƅ4*`(Z%���HC�3i.��jU��T����*�y�#,�+���]�u�`e@!bY���D\��9�v.��3E�9�8����; ���F�^Ei�������	P0������Ɛԝv�S&_Q�0�$Xe�0�)`�]���G�����������e8���n�9���t"�X,����	�Y�����,jU�1��-�i�FOUU����{��u�e�R }	�Y�k�4�7cm��*���xPmh����M ��	p��m�v1=�V�Q�^=z�ށ ��~����;tT�x/ꗣ"��An�q�Jnx_�`��Fi���q�g����{��y�z�C𘥌>��-I�f֘����]�%Ao���ȅF���!oaQȁA'BW ꒖iD�:����F]��O� Ģ),��B�>Ǜ��U�2vŐK���8�?�����a^�j����Q^�KHL�&<�%m�����y��o�<��<��r�6�@W ��$�h��������g� ��V�!�;�(��F�z��W����o�����C#h�!�v{[��dzk��
:�G?�
�Х��5ȄH��}
R@,�v��
P=C�:�m+�eIO�P�	�蛝����\�I�Q�H ]J��z䢐�����oNA���&ї��r�K"7�y�.�� �.j��~�Π�'���˥�J��Z�)%q����X�
���K�O�����f��pK�ˀ����>m�����eg��K�9�fi�����V�����b�dЭGlvot�-�d�k�Q�Y���R����u�]�������B˷d{j�$�c4��$9�H�>�I�V����d�!&@�2,H)�P�箊���/�Z��8ɃS7���.�]��������qoq8d:�S��b0#e' �+���P���#�;o�)E��r��OQ�#tq�@+8S�E0���/(1�	{�7tpr�05��s;PWh��9��'�"��"���7�6�;ՅD�2�,N� �i�)���~}��/�%j�[�:shT�ӗ���UP=��T`�H�_rT�)~������NC��a�����HG�<�a���T��LWP/\Tp���']�9΂[��G����� @�JEp�_�N��.�5˥F%7�oL��6ɤ��1�5u�L��}�=�e	��k��0)=U���w�`�[-Z�=r!�]�\�%-��:BN(��(�Ȱ�lA��bk ���{�̬�^���*8�c{�%H3���b�_ȶɄ=�xL�%�`/��8�qI��H����V�
`�oǗ���|��fp�U?%X�eo���T������/Ph�G@�.1T�ˢ
9g�'+��m�L��/7��ސ�K���9Î経 X�K4�9��ʦ�t溨.��i䱋0�x�H��yt�L9�y�z
n��	��S����g�I�ӊ@�k�B��<�S<5��j8��3v��[�*u���jD�BNy���=kjO�R�jd$xlw1I1e�����1�s������D����gs=�N�ME����
�Ly��>KM	�<�?b!py�z��?Z�:�c#��������2��� ,x���� 3��=�V��^D�ۣ�9Ӎ���׼"�]�3c	_������U<!q ���g�ۗ�>\��m6N���oyp9�
)b���W�xT�}��>��%^2+��P�3޳�L����z�=��M�|�ǵ=�-�]�,�����	