XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��I��f)@Ե�����j/ÃX�;P��%@�.q������֒j�mHlr���A�n�!=%:@�cT�bMiK��N��K@᎘6��T�t�g���~_S�R�}�l.�*QW�ZQs��У��f 1Μ˒�a5G��"�&�|��v<��2�qy�n���!�x�����Ɉ���R����n\���le��r�����v/Z1I��"����l p`M6L���WY~��
 �A,���y&�����p1����m�A�BC�a�S��"�QyY�����/~���Ӈ�I{P%��'��|۱ �2�#�����+3�Ԡ=q%������Ə/��)r�{%�ԓEq�Jŝ�[�Ъ3b3��F����m���A�A��vv�Ӄ�(�m��p��"R�|r�1]���m����@gΧ����E��f.{X�+�%}��G��NE�`I�������Z���a���0�B]9�D���H.L��lѰ[rܵ�ۅ���5�)#8����4�Q��Q9��UdTG��|��Fb��	eYay���3��'�/�@.ҳq��
����Q���S�Y89��V��C�\�H�ǋ$� �����Ca�KA�B�}���	��ߛ;����Z3$]�n�l ���-�A��4�����jQΌ$�5�mlv���c%��Qt��޺'[���|�������y�oE"x|�d^�K���>���[���ȓ	v�,��j����Cc��l�3 
���lr`��XlxVHYEB    fa00    2800��v��#��a��y�Q�tN8�{d=Zң�|��sC#���l����rha���ږ�7�0݉2ˬOa�*�ksn��Еޅq�p�re�+��$�����"�NL_�V�H	X��5J/{�B?#�<ѷ��#�G��ȄdpЖl=4qS%�g�,��vC��޵Yɀ>�EX��׆�~�����l��>�~�t�n�$P��DC�1]�\-yZ+�5t���f���^o��-��X�.��
�G���e�Y%Hv�(�
�o�7mS^γ� ݴ]#XN������'k�\^Kz�h�j�����
�*�i	L�Y��p�@���n8ʾ����қ���i�E�Ce���p���s���r��yU�!9�Fb#�b�3z0'a�!t-oFe[�!v�5\��l>4��Iϱ��Ux�:c�sduHRa���-�Mg1B�?ڌ��ó<Z��}d�~���}g1{sK7S����v#��c��2��/;Rh���*�\��4x���4�`X�P@���uSǷ�	��T2�	�e�D _���G8�#�M��F�d]�q:7d�FC��=��!!!�팒K�`.�&7ۻg� '��{3�ɪ�'��=���C�6���X�S�i�s�ՄX#H�_S�5��Om��d�������i6����#ЦB�	dr;�>���5�����e��e�K]� ?/�tV�m�"��,��2����i�s�<$7���o��b4KOVd	˧e:���C����1���S�$�fm���0V�EwH���<J�MC\Z�7��r�H��9�p8�䊲U.tT��7��@ݗ�2�V�w�q���y��965���#��<v�u���I�1W�v�0z+��M\�p���m��]u��lX����R�f����+i>.z�2|��j����:�>ES�G^�<�+4��y���x�PWx���ƽyd��an�lc��ZdL,���34����g��@��΃���M'��⮆�z�����1����[*��Ώ�^3�BPp��d�L�6�_�o��Qd�(���®�)B$��4��ư;�t�^�c�w)j29j2���ip���r�5������^�+��T#���)�B�b4���?�U���Q��f�߼z���i:͟�pŏ�Y*+@�hj}��]�kCɼY����7j�<oE�����k����&��9���h���ǒ�v}��Q4�h�Ș�1����X4��lJ�/��
-e*m�&0�$5]P�E�̠��&e3u�RHɭӹ$�o17��n[����@�/k;�����a[j�>��0/�xA,(�Y�zb���H��6�w�VR7ɠb0�r��YAr�[��J'i�O�Okcj�u�s�E��ƫ<�P��	����d�Sv3[h������,����wu�4��^���λ��.% �z�l]u�����(=)�����'���;!��[��/?9ѻ�ˤ��v�%�u-^��4�,l�Y?� 0����t$@�"��[��FP�=,�읡�U�y�o�îØXD}r-����8a�N�]�K��vB_����%���2�	�T뱔�����m�)>����C3���.�Fk�S��"; Xe��]�8[����Dxb)�$��=���ݻ�\��Q��1��g��_(q}��A�I�tiM���J�~3
���I�:vr:������Z�W	�Yoϱ؁+��b� o� �mn�d�}�i/"�n�^��\仈
�ָ<���b =G����dy߾A"��<P �賝�="��s�)C��f�ƆQ=�$����,�ޔ(�Qi3t�аz���ݨi�EL�����Dl�vp=��	A����j
���[�`t]r��;�^��{y�d�j�N�9*E"q�E��9�&���`��<]�@:�/�t:�?���fq/,�I�1�K+��E{��ބ�'��T�|��*�H��z"Ag'5sV��9˹�z�z��pY��lI�3({�Zxx����m.��gպ(~�^���9�ˡ{5mVP6$�89o����*�7��|?Ј*,�[��}�Z��yWĶ�0���L���)�����j�Zi�2�M��1�-U� �>&F�8l�*���A�$�Y��'R�0/TG7�R���ω�L"�]��R���g:2���ȷW��R&.-,2���G����:bX�Z��ޯR&�\�Y6�Da��(��/�k�1ۆ�Z�F�l��k�d��m�Dy���M���+��������8/�!��e��j�����m��`�Q���	琿Q�R�|���� ڕ]��H�ִ�IN+S��V�7��B�����zW�|�4�{����k�W��xWw9�р hy܌�_n*oB �e�_DM~9���u�̌7.Όƈ���M�`Q��Ƭ�*C@�ج��X�_����&��Y#K9��d�Һ{�#�7���q�G��egh6��}6�S��E[�}�B���~0�YH�� ��% >-���"}R~bε��>�񄜯���$����ķ��$�.�㇦��;�C��h$��.n<a��E�l��ن��&i��������r����N���t�k�Q�(�eD�)e��Ǚp@�"�۩�sJ��QV����+��㐏�}���P�v֦��"�XS�l��:�gB��ߪ�
'�j�$���9������#;T񴕾�6,f;ryqH�����s]�VF�z�r#%V�t�|��V�u�?4�Y��!� ���-8"��|2Ǡ�ef�1H��N&$�ֻ"jS��e��rf��7�(�fȟk�AV�7��A��xQ�����l>C���~r�h&�p�p9��wĻ�&~��SP�w��]T�|VD{|���,����.�ҟ������-5�˓�ˮmmv�#�:��tށ�N��0�{ED��vZ�]���)���X�Eh_�������1�*'ͱwv �'[;;��&#`�	[�����,��^s�'��o�{;���4h,`P�ɂ�`�����M�NU��|����N�J> ��s=�90!����-?}�.������6���rހt�ٱ���Ү[����>�����hK3o����q��GEY���n5-l��y"���E~�
��9�\�[x�986�N*�<P�5�@�.�]�죍��ݡ���܋,�2�k�)`�|��Kb�T����ʮ�Ol��J7<L�ӀCSl������A�C~�vV%!�KZ)At�C�;E+[�a���:V����>��U�%+�D�)��cH>c~����Ή&���n��k��@��`'�o�]�-F�ԯbi@����BOc)b	Z��ӎ���u�4>��x��V��fu�6c�'�����{r��}���;�J�x��%�綨���i�R�a�u�^��D��k����`���i�.�?U�#2[���'@�e����W��_��/)��oT[H�6�7�����r��'�F������a����`TT��$�s�\�ƒ\�A��8\@�/�-o_�Vq��4��F�se<G�~�3A���H�[{rh
�tK���Cj��_��`�dH:2��=���s���M@pf���K�0U%����]߱rg)>�x�k�:�2S�Ʈx��&�
�S`�l䝬����L�3sE�B���D��9��!�e��⺙�h����٠W��#8�/�F»W��V��L�Ugz5����M�����?�N��i�J�L����;�k�ML�Q�%颛�ьET"�qq._�#���y�lإ"@��=��!�3A�y�CӒW�ꆥN7��/�͉C��#A8�ށ�Y��g�0w1sBoq�.>��Kp$� ˹p����&§K����}�=��q-��yÂL����� ��ts\�-8�5t��8"�/=���ձ��FݣZ�����Dk$W���¸:�X�`�居�����藝KZ�%-(�����вѯ����˩� v)�ׯ�>��C_��s^���"��N
}:?˴�K����[/2tg�o;��G���������B�����Nm���]����Y��sfu�j��%�w2�Ջ�;���'�Zj��<x�hcˊ"� 13+nz�qud�鍥�d}�n���i���h��޴8bB�	}��@\!��H�\��5yD��hn#��l�J�o�0Y��o⫪jJH�����]1!r�X%V�Sȳ�Y\�&�%�l�(��aQ�n!�?S{_��B��	
1f����׼�ތ}l�*���P�vǵ��9��UN�	-.�\E�ZRWt����f��L�i{���:��$�^�^<�,�B�d�8�.v�l��-w�z�pW��g�z�_�Nos$��}� j�PL^"6(3��u��8X��3tJ<4Moy �$��s��}Z�����җZ�kG�f�,l-&���l)4hU��~����21͗�]��&�����眉ӻͦ��Gaf����Im^Е�:ӛh,Q�j�9Z��&��O�<���y>W ?�*h��T$���nix����r!��A
�al�{���x����0���6���u|h�be&.3yp��Av�q�^��r��G%"Zi������p�]Gn�DteH\E�o�tYm�ã��.����/�yT�1��:z�嫣KP�zA&��t*'��i-3��;�t#��e�@_�')�_�B�Ӝx�|�sg�(��T3�VPs�lgDX���nV�<���|Y����ۋ�vY5/�E�`��ٹ�9���*+���K˴��%kF;w�3$��R�+�c�ϖ׎ޡ�>���d�����!�p8{"k�)rG�\�?���7�J���)tp|ۭc
cq�;�:���u}s�'�b8��](��h�F5�d}ƶJ#��b��g�� ��6�f�r�Y�F"	2���S�3���<����O�����<v�H��{P��5���e������`��ж_���CK��K� �	5�[���뇤�({� l��C8bM��V���L#���?��5Ύ/�5�I�D����e����[J���h%odκa'x�g]0��m��t�-U}
eIe�B�}���0x��ի�E9��j���b��UF��3������!�v�����WC��ń��,�qs��;^I#�E{T����	����ky�\��j��hgͨ�d���I�{VF%�~c��޹�o�I����6e�Uʐr�m5��A��4������W�h��_�N�7�]VV�5 [h��t*�t!g*QNݬ%�ۗ�Udq��G��^�8��W-�̵0>�D�=��a'���%|�$֗�[�`2���^|I^�������gA���55���M1���ڀτ7�%�*8tN�/[(}�n��� �ޑ��X��Bb)�2��@|�Q�h���ٯ�?���. >��aC�I�ND�Ѧ�?aÉ����p`�^�D���
`�`�#L�{C��C ��`P�վ�*�+ț���:��)`Q�oO~&>^��P yj��&�ӄ��#b��Ȝ��8k#�h�C{���O(�@�,��;�PI����[T��Æ��lU���`o�S�2����m]ZSJI�O�42'g@�C�>7�n&WJŧ:;��i��#� �ë"�26�x�z�{����i[<��斶�A���gК>1��	�~>���9���R���GZ���:j���z�LO1s�KP��[4�`�O7��ݫ�Vl��"�\lI�Y�~�6'~�n4
���C����B�.4m��Y`�����#�\.�]s�' �^3;�L1Č�(�����r���/��
k���9�^�\m���b.b��>��U;���.��{c�Ւ��/��;����3m^����-����}kf��pO��Ը{��(�9��6�p{g���Bօ�u�g` ��~��6�*p�"M�u}�mǥ�����k�s�'>���p�Y����;Ϳ��Z]������m R��bO���Q1��+`~����ފ�L���Op�͑�JlT�ho�������"4��E�Џ�rMv�#E'�� a"�a�$:՝�y�:��rd�����X^���1��[����Ǩ3k� c�Z(+X�sT��!���*VA�[�4@�������D(}��	*?�J\8[Z|(�
�ОXg��:�vg��^s�d'p�)�&	��a��&�cG�Ǜ��`)c;ym�d�;6\R�3
��ZX����H�0�RJ�=����w�͵�QxI�7	=}����aSC����x��4+���/�C��>�q{6�x�k��w�Ww�A�E�e��5�H�@#�RF$�t+��'ŭ@F\���� ��|�c�x=LOJrk�
?��3�d���?�������=�
6�{9��CK�J�W@��Nrc��j��	�\-�@R����ష�-޷��>�'����YrNfl��K�J�/�pkmL׬��2Jwo�љEc�H�a9���j9Kr��~��� �/$
B	G����F�����q��2� @������.-8��YX�Vb�ݿ�&T�M�z��h�����,,oΗ9]�i�s\7q��d��&�p�w7\X
�~�ē9�~{�$����5�R��P3$"W�k5�M<8?^hFF��()/:�x��Κ��� c�|�����}�o��RU���Z��u��os.�$���:���z�廟h����6��Q�6L&���K�uHGjQ���6n�K ������U,�����絆��U�#�S�D����ah?Vչ��H
4�V  � ���;�AK���F[�3l�e�5��m3Ѳ����@v�4���]s���8�^�g�����fU�^vū.�6��T�{a'sЅ%}:_}f�V@��tfC�hX���*a�q�޸Rܿ;?��	��jK�	uV�P��IT.
Pj%Ozx���-"����QҼ>x�
p���:#�)QԜ7�8XJ�
vZC��r���6���Ғ�Q���	k�-�6�v�����p��#ԗ&T��³�Ӫ%�	�$�EI������!X�8� !fx5���xz/),��`���X��k�E+z����	^�R�LnZ�����ӑ��J��
cJFL��� {�b�]ch��T��V�m��6��weM���4�P����=?��5zf�y�i���z��M�&'w	��iA��l��\�
n�9C,�l`�Z��0dF�	�u�(��7�����IP�^��!��i�
�pRJ���v���C�jn��ԆȮM�xr4�^�̡����h/�����=5:��)^�=S�����m�!�@�H��M�n|���ը�< ՙ����S}F��g��C�sg���;��^�M��cO��6�u+
EVl��R�t;�<�������X��� uX�xُ���z��Z�M�Z�3&��T
>z�N}r͗5Xv�c+~z��a�E�,�ʹ���h�[G��c�a��0�������sqc���P���˝�Z��/V`��Y,����AN�h}��"�`����q�5��N�E���>o��a��Z�A��8{_��z!�kHh�h��L'�5��ZQq���-����^���(?f�[~r[& K/+�또���T��w�Y�t�#�7ڛ�,���w�N0�p�3���;`�`��~�����ǒ�*0hA�{�C�3j�(�^�B�ki�]�XFa���9�)��؁�gƂ<�q��&���/g�B��q>@� �'+�#C�4�y��sثb����%	��M�ix=��5�$�70.Zq"w����������JI^ 	�����F�MS:j&)�2��8�i�x�'�UG�{Y����W�w]�䢊۝GuzNc�.Q�k�|e�~Cs��mo$�s�.9R��$��)p�t~a��?�Xk3��G*j�]�l�����Ks��ɬ�R���*��M�v\�x3��p�Q|R&�z,Y��4@�B�X�]�h2���Y��΋��N<g�vļ���R���1�^�+J�#��7�5*�>���hG%�E��7].,����	D'��1'd�%���M�Ф�nd1JX�8P��k'�`"]P�T޻[��|k�aݙ�����cnJhu�}��oz��D:�{"3[�*�'{H:s>��m§�q��lΰ+ʋ�ݚ}%��i�>�6��mvh��䏩�v� ����I�_�p~�(�o��{PY���Y6g�k^�_<!�o%�a��:[_��%>J� vu:E�E�g�CD�q�2�T��!��
��v�t�kn\��\������4��*���wlm.{S�x\��,j;݊�>&;6l�m�bZ.�'�6!�L�F�6}��� ªӿP���G@ұ�0e|�5b��jljp�[W5�͘·X3��Q���A�����k�|��g�uphy�ŉ�C�Z�}� d'�|�����Z'�=ʌJ��j/�"g6��rC�)۱�	Qgm�q�E��R���u����'� �6�U��Y�\�}b4l����e���Y'X������P�vQ0L�}g�9�hT��%�=�R7����P�4�`/ԅ{݈K]o���G��p\�������G�%8{G�[u���p>Qe��ru�аW.�����"k���='SE@�q
bxp��j��W�u����?������D�E����Yĳ+�
<�=�W�)uk��UF�./�]t���w��WR���jZ�j��J�,Ė���X��+?�)�'Cz�6Fj��*�mut�VyU���F��H\d����!'��I���x��S�����B��V#E�Ux�ن3z�-:3[)G��"�$��xg�=E{�py�7��/c>��uGK����B�>�Or[����1��o��mI�� �bʥ)
L�΁IV]��Ǌ��a%Zn���撊�<�-Yi�NH2R����D|&On_��_^����k�u۬��2�Z�{7�H��!���@�Pݻ�24UI�ԝx�=K�� �����)I�ڽo��ok ����]�|�U��S��@=����y�'V�����Q�	��>��cVM H�T`�1������M��D�;�|+�sR/Ὢ��<$�ސ�2�02�>�\��p�g�'�
�5SZX`y�m��]�>(�&�K�1@#ܿ����~J���t֌�����P-u:�}�> f���t�
SA�=`1|0'՘h����y@�a�R�-ƧͲ>� T�n�12қ�M���C޿�����M=?V4��Fc����� �JL�7�Ъ_�����f�e�%<��P��z�xk�0�u*tIng�eL�I�s��@���ܧ����	X(���!F>�o�ie�R������1ш�Wr�$g�>q�3o%Ypm�n�Rk�EC��(�B�[��s�?��
o�)��py\/j�]�0�L׏z�( qqfI�cZg;MԠ\|�/iz`r.% v5�"[�צh��d�{S�Q� �lu�c�֮��L|����g��{��|��i�2��mG�>e�X��ke�U�H���\�QR��z��'�Eg�?ŷQ�=�~�O��
�o��nO{i���f#���.���Te�+�"���H�#�zO�.��B��!����}�t�75�8�XD�;U���[�;�VU6Ɵ�T[^��'�>��!>����C���+�=�����s�F����I x�#�h7	O�]�M���qb _t�p�;��b�3m�ᩴY@ֺ��;9���Vw�+�Xn���N{$��U�96���j�̧�'<�y��S�A���4�h�jP�E��.W%HEv ypi�㶇��A���`��5d���$�$�c���za,�TYxXq�k��rѿ;EI���jl
���r뱳�yʷ߉\vq���=�]"n��ze��|��m��nj2Z�{�t�+��$Hk	��j1Q�6�B�!<nhƋQ�4 ��*`h�!R��<�ƻ���������g���A�"�&	�����m�:;�]18l�<�4�Ǘe�&l��?����T�Þ6�CC>��p\D˴:��:��8���y��Q��0\,K*uH�#z���NzXu�	�H(�e��Ua�m�$i/2't@�g#9��H��8���}C_M%�:v��C��r^OD��;0%�w��E~te=?�:����XlxVHYEB    5ef5     b50�-���,P����k ��Ao��a��,b�p��������+x\����a>�4d���DV��Ҳ�����
az}P~H���6���/�4�) ��(��DC� it��@�d�q�>�n�8s_��9<�?�d��U1�-��y�&���(�LO[<1)�Ԕ�=q��0E�	�z��	]L_'���~������~��q��������ζ��<=�D����NJ2p�
�V=ʪ���3+0�8evvMARN8w�S�E��yF��w� ])�H����n��[��xb�<_��s:����؈~4��[˷Bm��J %H^����xn����O�NU��vꈏ�T.A'��ZE�PG�ʂtˏ&J������Ά�������A���z����=i��li��^�	</��`�A�)Ѻ/m��PMe>8��S�������<�v^��D#S7�\��&~��&��"\`�P�7��Cǰ�ܽ�*�Z��	��	��6�]���C��FЫ�)'��u����u!��>p<��R���IJh=�7����+����f����U�r-�sy#����G��"Y��fqf�%�z&�J���?k��ύw4/�xf�Q1E'j��NW�+�p���>T�̀��%�q�M����0�BEs6�	���!ܼ�J\��c�5��^pQ����|�<�t���	���D��	Sn£�;SX�{�W˗Y�)�Qg�l<DA���(.Z2�W��l(��J��T��K�o���58WC�7@��
�MC�p
tTD�A^���S��}��1q�:}�[�-�Ű8��2\��Q�)��<Ir]��a �fI�}aC����{b�V�]�Ѧ�hI���z����+R�A����mB0,��[��h���v��&����)�t3�!gTfn�Q��!I|��r�m�<�-/�����`E@�[C��Q��Հ�2|f���4}c[C�xj�`�ro�B��8���)���=��nˌ(�Ђ�5T�&������+��MW�@�ͮ�p�!V��j����~��pRy/�Wx/�#l�sVe��E顛�E`��66���/gęM7�	J�P�U�`��ZtFtS��G�т�h������hɾ`��6G�gX��=�
qx�;���'�Z�X�mfu�@��Эr��*��i�$��+)�^�PNOP�\�m^��h3#�YI�\  .aU	;We� 
�6�I�Pr���5g2�8�)�R�v0�b2��R���l"��%auq����0�ϖ�C��ѩ@X�.a>|B/���g0��7�]�%<g^9_5��u���Nnl[񗄉u��qwO׵:��n�y��_-ώ�Z���ORO�%�JƔ�_�]�D�@��:�
S]���S�k^_��ަ��fx�δ�o���F�pV�q�a�\٘7�.M�8�@��=�8���J ���z�T�Xn�#�k=C�w�c���2�/�{k*X�x��f4�kXS��
),���E�����|�p�V�^M
~LY'u�]�f[�}pl{Q&("M6?�� pF6�|{�g~Df��^(H�mr*٘B[��H�0�o���q�~��La�N���о0�4D�:Oٴ����q� �R(3�08�I.��4A%��BF`�
YqB�,��ʃ�X@ܭ>��6�K�8�����F��\8���ϟ:O�b��gփl!�Q9$<4�hSG�*�/�,^|y�����*H�Ty/� UT�H�b(�U�C��"�T�\��)��,7N�BFL~�[�����.���1���AO��E��+�@�chz�[h�x4�c�&�y�`�)�n�J�ë�rh"�\%������}�b<�X_������ml�0t���+Q�l��ܩ/�6M�@�_q1���A�	�)OM��:s�T͠)io7~U2�Ap�����V!m7<�C�3f.�I�q�T�vO6
����|z��$���f��f�	wB����iU�9�$��aZ�\e�/2>���{y?�TF i7��"���ն�BjO[�JC���G�����N�|�t���iƀ�L�n7�y�𽴿�W����P+�ח�����n����]����2N���2��B����؅@Ͼ^_�N�v�Tb��|?�ax`�G��m�"j$�o�����%3�,-a�0�u��]�E[mT�7�]H���n��ޛn+��x���5��$���da�)
 �"��,���sbh��@q��n��]�p|�m�$�l�E��i���21TO�}�����z ��w��K�|�C	�W��NS��2���m����ܗbְ�?ϒ����ſ�>��fr&�sբ܅��_F�y�� @s����Yy���'Q��F�߳�7�jFI*�(���v-2�G.����'䃧v��G��|9��I��'<h�&)���q�ȃ�.Ż,H���=h�g� ��i��|�MG�6SldU�K�������>í^&�};��'%my��g+�Jn����p75F�ܷ�A0p�I��s"�)8#ȴ34�LZ��M���	)�N����C^6��v��xu���>nJ�D��I�b������9C����L�p
?R#��E GU����5w�'�W�����(��}��_讏ă��� &tk�TC��@80�C=�˶z$$+�(͝��SP֋���L2uA��f��0�el<vs��z�P�����Q��0�!n닎����^��d;f�:s�{�5�YV�����~j錐<�)�#S�� ��߮�a�������2+�\w��n�7M�!�5mƿfؖ^��qc�|V�����nB�I�e���