XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��b�d�$⭗ZU��e7;��@u�:�wn^�fL�{�D(0�a�n�"٫]���c�����ҟ߿�Ђ�H��V�%ִ �ΎMvG��SN����3�P|9��P�Н�gj����}�W� .`y%aC��8�)H��E~����@��#>W�A���tO\:����e��[�1�)��΄$�ei�ď9"�_V+8I���s��ip2U�W�S�Y�P�v��p૨�x�w|��s��-P��hLK��>�B�ӵZ>D��J>��`MF��ynBR!n-v��ޓ�nNi��=yL�i��޻�	��8�@�k��sm~u�6��=�������	�h��;x�;B��4I��- ��a�MV��j�b�%�����ԍ̀i.����hJ8r�4��=4���+Y�,��
��̤�ׂş�����A�� ����~y�H��b�]��5�7��*s�t]���*��H�Y/����)�/�Y����3�������St������e�{08���"/�����7;!��\��."���&� )�\j���6�f�����`�NaI�����e�Z=���y�||6亀�05����+F̧4؊�nY���3�����췸^8cǯSeOW�#]�5�B�a�חqz����qI&G��|����[�3���&��A�42��?K[�Z��	�Pu�6�C���yK����i�f��e�/!���I����n�<r��|���D��`�.��a�W�ֈ�T �FNXlxVHYEB    2fbb     bd0g����<L
�L�$)
���C�}����}�`���7��D^/<�=���sJ+�i�o��Ui7TO)����̖�a��Hp� .�?�%Y��O�",��S���5���eZ����x�U�d�D�K�l���281Sn}ʯ`������ƕ^VW�?�F����X3�T�:��() 7h��D��M6��μ�3	*f/�>l�n��fj7�0�Z[�vm=Xl&Pѐ��vC��~�uG�V�2�p��܃����b[\3�zO�	i�%dt��(��p��G!T�uE}�Y(l��ӊ�7.��Ÿy�p�>(�4��Ԑ1��ol(1�X���K]�׶�&q����a��j�{>�/2�ŝ+�mu�p��j��N^���{�Ԩ��͗�������}��UA�_�����E}�����!��%�M��q����񮄊�!��}���B���&�h��%er��s�#,����%*�e��L}B�k>m�'�BL;�&����Q,O���e��{v�� ��i`�ƾ����D���JΔl�/�������9P׽�-*2=I�~���;u���e�$lR&,'���z��o�]����A7���
@�I��Y�A���˘�0��J����\�DY�GjK�h^�
�쀫=h?^��tc\�r�剴�}�x�ʞ7��ٜ]S�w�Bw6��0OF2G�W6�c�f�&p�`��_a�k,������H/��u�]�b����za�p��9�� ���13�Wڒ�݂c8^�����K�/4G�4�\ԭ�g!�Ӣ=��S�,��'�U�F�P6�&�%�*D�.�m�a��!���S�g��&1;ƨv/��PӅ�Ch�X���pttgqT+�o��b�$�X�@c�sLL��hX6 �F=b�҈XQobp�37�&�-�p���V��k����ld��%��'-L��ڳ)�7�nJx!����0ҁ��*Qt@n���[�y�?�C���+��~�3�B�@H�+�Ex���f]�I����ܞ �('�ɡ�����W��ðK�ǽ�z�~��/���T��W�c�経�bN�v�/�䱎Z���HS�
fT?ڧ���y��[��6T<U߀��~'ʓq�����A�)��S��peaSu�%��u[�dj@V���ƕl6�e[fn|���c&��Yl���5���
bM�z���D��l*Tb����n���#yv]֞�X�=K��N�M�����#��\�p_��~\
��p��e^�)cㄷ�6�w�U��K%'G�-eGwFhŁ�Sp��n����Qk����Zg�
�Jf�K�o�=T����ӯ��l��)�r�Z�;N�@"��/X��;��	I��2��{�Hj��Q �����z�L*#P���I_�HE�x����߂�]Ø�����.ּ��km���J�;�&�����D��I?�-��Ӥ�ՠ8nc�"E*�	��z��ө�׋e}��n ���L��;D��j5b[��J��\�'�Λ,.�t|G6Ux>|\��0����mRݚ��㮮O�Yi�}(ehq>T�MÉ]v�@M6�{�|�R��G.G^�c��{��7h��<��<J�̙� �0���L�u�����v�@��Q� �ک�o.�߽|�A��2�ݮ"eJ����m�� ��ә��eV����ߗ<�@��c���4E����]|�@�����P�or��>�G�Y���������2#��,��M����l-e�PޝX�j�\[�\�X����ȣ`R�sp��By�%��> Tr���_��Q=���ІϏ�c#ê�) �.�_N-H�{qN<` Pd^�0�=��'�Fx�d+���u}�`i0R:T���9��)u���+����7_�؊�.�OP\��6������3��=�?�����o���m��!�$s��+�:���Q�B�?ɨ��q�xA���H_Drq�`nc�q��|�gWjE�sS��.�Xt4���q�q�Iڝ�3aiF�ɪw�?k%pN(�my4��Ւc[�����g)!?��p���k9�%�	\X$̾�)~�v|�*����(U��[����4���?������j-o�.�n����6<��y�kB����׼;z�tZ��B�ZZ��^1]@�+A��^�y�c����˟O�M|�k֞~�*����Vz@w߀h�Mrl�
{�$#	H��b!iV͜8QA���{��)����{u�
��ְvUR�/%� ]�"��}��9簐J'cx��,a0.�{��ۭ����iw:#���瘂����,V0�{�gF��>��5����S��*�!|{��^w�dVn��f$���ޙXv�����P"����J�[D5W%VJ�H����JqYx4nq隗��a�>���5~��tH�K>�'B�p���!�c�eNs�@�W��F��'F�3�	G\�|��׈"vq�>���oR�A�6@�4�|I� �������2����!��`�N�U�uQ=P�i<�qv�o�3"��􄼎�$��Q?ѹS�P /��*C��z��Z�5���CGm2��Y�+�^
��<4dnd����4a��~k+��&N���4�U�On�(�]�Y��	+kB�U���3�l���zD K�@�/3��G[[�"�5Ӻ�ݹ�:=D�6e�3J�&��8���$�����;Y�L��ڇ���E{��ib�m�&��!�y�d�Z�	�h�0�i�[��X�*@tqn��#�{�(��~�i��`�9�x^@e������� �n�_��Y�Y�XYl(#�y��o��_%�JZ�!�z��N>�24��ApS�,�
hG(�엘�Y�
*�d��������ˑ��5M���tt�1-��;ܩuz�y7�2���L�`��T��� �_{�c�9.��y%�`K���+|_�e"�l߮&�@���PzN�u�Ì_,��*Tj�'v���$Ɋ-y�V�OUe4���t�́�>j4E���&J8_�Ld��>wc8� �������b^�Ģ���a'w�