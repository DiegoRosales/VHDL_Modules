XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��`l�g	����A����}k�����OF+C^6;�Ծ%w��T0���o^ԟ�+�	�P��@���Ł��'7x�ؤ]�o4!�9*=n�)����]���4�����d�;jt��j/*�CX���l�B��)�9l�
�/��؅����:�=�H��^���.h!�5P�ƍ+@��]tа���0�E�\�6�^��U"����:���;&5�}Z���$��gk�&ĝ���\�#4{��3��5�hL�N>u�{}kr��Q)��6��%8~����	B�p�r�S�9	�$���� ��*�U���P�N��Gbސ��E�0d��s2�&g�H�Se�*�d�)��ŵ��b.4[�Ӑ}nt]�q�g��9t�3���b^.���y]ƣW3����r���c��O����lc��%䞮��e�~=�c�ħ{>DI��-y�%�O?�����_r�+1��+��H�{��G��������{::6�a��A��>���Z��Y"����J�M�+atٴ<��!�N��i�;����ϱ	Z���FB��w ���OڣK�ʖX{�H@�I��-�Q$�^.L�,�5��`@jɰz���v�7��/Y�PO`'��hƍ����w��Ip�))�T��a�!W�ыN�㘵ݨ��m�y������9@z�e���,�PP�	��Cg��T��Tȗ�A�HP:<bvPG �Lv�����?0W�9�b�3���݅U��]4�}�y8}TV����J�l�e}�� T�����#3���XlxVHYEB    13ec     7a0�0qP3�03���Ҥ��W�$�����F�2LP�Xd�Tq�a�4+�a�3{gxOX�Rb:yz�5h���Y'��7���v7��U�g*X	)�U�t�m<R��?V��>��T��(����Ĉ2�9|�UG�a�&�i�%9�Ռ���-"r�t����W�1�s��pGͬ�8r��� J�%8�4p�Q����8�� j8��-�@Ei�}����|Kډ6s���wwd�6)�$���l&Ĥ��@��ҭ�h��mC���gV���"���]��Y�X_����˻����"���|ƽfPc�n��S��	�N����x�F�-Y �/�p,���9��%ୈ਍	5O��R�%�(���nvs�~��Z^�: /fK���*���(�"q\F��&�tL����4V}�& ��o7��ο�4�L+��\��N�~�S����*���?|F�	2:?omZ������a�%ZЄ5�awG<��V�m���Ed�\��R��B�;�p�\�E���5O�"��[)�S�53�]�@ܨt������0s�f�+���F�|���Ass��Ö��.�������&��֗���]٧K��;	�\���>��ȫ�ܙ2#���8.
JA.�k�@r���
��#����x��**sa�~�*��jh�mB�f���4$̔d�\F�ow��Ț
�l�k�l������k�7{Z4��FqPy����@���>�8����v�V��M��&LH�j:hfRr:���x�Tl7��j�ԃ�ܱ	�[�N`�e���M�è=s�Y�!iq�س�H		T��h���h���Z �\]+f�Tl+y��_��������@�R-�q�t�Q��u��LpC����A�VvϏՊi�3t���~�~ȕ����=#g��W'�� �Xk0�a�j��"I�_��|lv{�:�������A&'!}��mX�;�9�li-�L��R���bѵ��2�?5o�? �k�h��I"�_;�<I�yZxi��Ŵ��Y8ox��h�T��z���3<꾤�̼��5����J�{?-�������z3e[;k��Q����HN���{���w�)	�ޝSG8 ��������<1cӆ�ȃ��W�)��j<	}�[{pa��sʃ�^�k�N���i<LXE���u���:�m2,T�����C�哺|���3L����g:g����"a:��B��dD�+�/�[��9���Տ�Pۻ�f�ߤ��Xi�A�1;��Sc��r6�1�:h�,x�d�y�q�Z� �r��(G�i�����r�1�di�M7���ǟ�<-�1�-i)��ㆸ�A	~�L�坺A�;�E�H���h�gGe�Bs�q����eR��ARYr�L�A %�,���I@�_7�wu��G�4�т`�3~��9p���j'T2Jk�k'�U�y5�����g��<(�:�j�m��s�{���uj��L�;D��pEt��5=�����T.`�j�t+r9�rUW܏'�N�7Y���^eo$�[9�D�)�g������U�ś��qq�4�e%�zD�ݔ�}����J���4�[�8m��!3�4�Gتe]y�c��8�
���8���|-/��On��D�17�E7��W��x���:-�W^�C��N]�w�����iaoM!������9Й'
��)8�@~<�P�]Q���i3���W]��W�sؤ�ͅ����^x���4��w�v0a��(7�-��In}�7ΐ��2MW���g��dx�W��"#x}�.�u<��ؙPףқc�;#nǶ�GSE�yM�ӹ���m��/�{оTql�)��j^j3�.p
3�RY����U�F���P��*�xJ�X���d�ж|�o=b��<���/��(��2�3�r7��_�������⭄l����Y�0�i#���u�{y׾ �