XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�����v]ް����ծ��j��$�vQs����k� ���&�������z
���M�.`��fq��PG���>tgSv����n� �Rȫ'��c-�F�5͚���s� c�ä3���R>a��׫*�TUV��P�5�94��}aB+D]3Tv0(�y�D)*�X�)Gr
��p8��ĸ���I�i�|��E֌�%(�F���v�\? �N����0+ZF�5�w���J�8�ﾊ`��8���>�Ww��B��ŰK	HIO͎�eGF����k���1���+
er#+���n��th�Q( Ey4����y��ֿ�@��'���ıYv�Ǩe|h'�g��W�O�Ӌ��d�h:Ώ<'W����,�N�w˼��bTm�d|gl�%Q����}�})�S�ї#
�*0X� �!ő�U����=uS)��hk!�O����_ۺ4��@�Qp��y)�U+�wKi�9��f�%D��C�����#ȈI�k;F�������Ҩ��������.4E��'Ye�Q9��Axtm��[]j��$)�6���~�����-��~��Yj�����y!Y�T�<�G�e�?m�-����Z���`�/��'���ozclϢwdEPJd8�@v�����-s������t%�~(1�i�\�
���S���d���Ao��rU]��Qr���2a����ʮOv�?������|�<���(�_
�$s��픇h:K)�B��\)���7�;�U����k,��rP�� Է�s�XlxVHYEB    1445     6e0��=7^D�$�X�כ�����G.++��@'9]�u�vw��A��ix˩&d�d�Fc)�}� \s��%�D^/fSb=nҪ�z� s���8�?�1��A�� {�,$)�����]$h6��Ru����b�f	:�=�i����	�&����Y69H5Set�RS�.�8���qmz�m��.O�Qz�iO���ĭ8��m�x�rA�q3����2�]�U�#��{,_"�5��D���L

��bg�=�,�u1����H%x���q1�4 �q�����&������ �������H@�����x	��7����҈2�uNciL�9�8�[k���%����3$wq��6S7�AeE�왒zL���׹3_�u��] �6
��ۼ5��v��SiK�,6��CF-�qQ���*x20"'I����/�1� H���N���G#;.�<Gɥ~~'��a�F� ��_^�h�7)��֟#C&L��ި�v��խ�]���oY�I�T"�-�\�cq�J\�,�<t��{�iB&�i52�T��nBa�r����5���r�r�Q�&V��bcl	�̕� �� �2kw�a��O�x/�WC�;TH��[]O5���k�
�����y��Z|�i2[7�7���%�7x*������ْ#2��ª�cz J���� �`�n=�`�\p��-�6I��tg�C�3(Y}c�i�h��3�P���0Y�J��v��"��i��h��T8|����fl#8~gQ���0�\��͚�n�M��v�^����F��sX8�UOFsfr� �Fc?x�c�
�w����V�B�=���Ļn���<C+��X�

1.3����A�-�Mu\���^��!T���x�ʨ&���P��M�j��}��x�<e����Ј<��Ϧ�w�����\��"}M�;�{� �G��̇�+#<����B�#��O�,Q���������(��҂��&/�`�2�"��E���KH�{��|��,p*�If��YM,
�	x{1��!E�r@R	䝨��6�����46a��I ��z���|���gNM�A��3ܸ@��x�
"B��L���B�yu�~3����� ��Fx-��H�ԧkψ����D�L=S�W��.�-�TԾ��aF����3�eu�C���V��5�0MH��i�k2%yAS6����U�xzK.�Ma5|��m���]z����<�M����*I����YE4&K��������չ��=di�@^0p�(���t�g[��p�])E<8��Ԡ�4���x���t,N�J.\y=F�z����ޱ��(|������7ufC��9Zz+A�g���O�aL��o��br>�|��FD���N�#�Wi^AG�W�9��;�o
歡hH���H��ϙ����J6���C��/v��zͫ'�l�7^��6={�󵝽~��r�nF���սnjqܰd�����gp��"��;���6��AЉױ����A���[=�=��G5oj�m�s-��8�-�`�P���0?�~ �T�$���5�'+�[0�^B�֠\W$2=���h؆��E��}�f���BM/��T��~�D�kp�Re"} �_�^#�p�uȆ��N�$ʧW�6����◉ң��7�'C��2�sĘ���]��=������>Z(� 6v���I������vл�3�59��R�}� ٗ���[L^^t
��	�P`�@ۦ3<l�?���+����w�