XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���"V�K}@��f�rB�J�5���<_@e9O���y��33(��`���Q�Y8TAlA'��,�N|)�M�ņy�s�؜}tyg��� n1���3qH�ě,E������ė���ޮ3 w�ۦ<��n�lE�]<�y�N�k"8��V���[�Xi$�������_�p���n��k|)��Y�itO\����s�R�ƈ@����k𓩓&����9��r�$�L�������υ9B�)+����� ��>o�L�������L�jm��'-������:����`�p5��m��Db����hxR��{���Yv�M�Q�������T��+[ Erz���%h�o����{�P�n�f � �r'�_.ތ�ey���)A?�xf�ܭ���35�rpk��ޯ1q0�-�.^�ʑ6"���V����Aa�g�@�3�6U�)P�?�[�R�l��!����20ob��� VІ|z�a��/�x\0ϕدc��\1�;�"�ߎ��*���&_�!ŬH	��I�1=)6�EK�����[��h &��hh��d���'�nEY��{��z�}��B�sDJBn~���Hk�dlJx�N\9-x�XUu	���)�,���X։┴��g�ןZ.yy�ͻ*m�g��.H���5�5�2'D��O�ev}�"+Mn&�q�
n;9d�<��%)�t�{[ d���*̃NAC0�1]�b�8dH˯F��i))�k6H����~��8$�*	�c�XlxVHYEB     e37     6d0�ŉ���c�c<5YӼ�ck�+��Y5��/�%��SO�˙YT�߾`��rM��G��������LLz|I��I��-�]>��S]����;�-��/
��1�����3��� s �673P\�L:��+m(�"j��ݔї��ԕ>$N�XsD>���ћ'q�Ҏ��:\hD/V$m�
<�[ʗLj9�7=p�A$�꫔�ʫEHꡆ��>��V�n�ͩRw��&��iy��� 	E���$|(�ȼ��Aw���i����A�#��zd��f=r��`/�K�P�������V¬�gӨ�2�̅> �>Dc���Z�lm>�L�nViϧ<�J�Ay�K֬m1(D�+P�����UX<�0]���o�<�2��M���`�j?d�3���Kۈ�t1�2�*l�����3��9��b�q��ۑ�W-L(`ZF��)~�|�8~��J�}�4�68���Ux5�S���Y���o1Ύ���N�e2y��w5~¼:�y�1vf�&I�B� ğ�P��͚'��6YX��!��b�!HL�@��e~@��i���(_�w�HǛ6���80�#?��.E�gp���f�|�(=7�?Z:[O��G�&7Xv����1��c<�n@R��^>�B�� 4Z����}�U�ð��V�����GN��VL���-����p3t���9�	?��O���+6mVdK0�J�*}M��ִL�D��k������ыHK����es��v�B?(��\�J~��!i����PQ�F�%9�ksǂξAAe�o�n�KݍkA�!���j��� F�޴��%Pp�!�x=�U�zmP�dm���e"Gh����|�/�B���$:X��%�<�u&5��������]��	����V�Д�D�I�1Bٛ�����T��^.k�͓�8VL(�|ômf��L_w�1,�<���֡����� ����u+٘��^���M�J����ƾ��L{f�;���_b�I��iS.Juz�v�So�(��wv�-6#����ǩ��NE��I����{�t�5J�܍G{L��jA�5r&��_�)�8q+i;�
E'�[�TkQhD�D���<ǽ`�^]�$��P-���<K�E��/�?����뛰i�j:���m-��Vg��f���1�_M�����~y��?�h���"�ZN5�Pp��X9y^Ed�۱�������4�g���)B��*"|mQ.�S;r+[�ƑH�P�W�����55�ܱ�ÎB�y�@5���U�ꤍ�l�	Bѱ���nDծ���޾<�z�,�&��zk��2�x�s�,/���Nu�����T�S�S"w���^���AX�C���0ۍn��X��W�9�xe�o�PƑW�{�Z�+��!n���Oh݂�66;l�Z���!����{���Fe�`���ox�pʚc~J��y���*�SMnǒ��H�Pv}�I9��w�ªD����	%!0l}{�|-��]�c��k��.����%YV+Y�P�f�t5[����*����!*4�U.^i�󐗮�KL-6U�A�Fmڪ��_�@7LN�LTF��a�*��|/7���.4�
�V�>U�@/�5�����_1=��.�����.X�a8�������rqjx&�e���6�ȅ�-�b�#�G �҉I�jP��Auɛ/���V�mu�K���2��������O��J�X�"����z�ѝ2����D6��ռ���9