XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��[��_Cy�����A���mF�f�ǄNIk�4{2x8.���u�,u
��)�)צg9!D���}�U�p5��0�g��;3Qy�sϐV��lP1�ǽM(�o�70�W����'oڐ��st�y��qu��^�\n�S�*<`o�Q�a�~� �#]W;u
��3�c[ r��������|��)� 
��fJ�z�[��[�"~�ci|��W&؝����6�7|�����C�H5 ��1;~��C0��|�3Y�h��/2 ���q'!hj������k�%�܋q�@�k�ƅڞ��d/+��@�4�]Uy�/�.e�^�`�na���h2��`���	����Y��H�E�7�̶g���3R�BY�`9�}S�9��}��%��Lƀ�}�B�08� ��(�B�v}D��]w��o�x��o�ths-}��lת6b��,��v����d��?eM��X�~i�?=MF�i_PD�,e��j��Koi�����B�S����t�Q�2�v"�n9�l�Bi6>��?��H�\��E���u<m�^�Ӌť�\ZP�6)>7`}���pXN���3hT�d�i�{�?�� 'Ә
�	N��`zޟ2JG�T6�;�#"G��R�g]k�[L��6���e��������z��K ���V~]��5��*�9�a6m����.]5��t{A�����Rp�{��NK�@�8�&Dj��O�G���qC�Ύ39��`;t��(��{2�k.�;��0��̴P�kt��ȯ���]XlxVHYEB    fa00    25b0��^imB}W��Ś4�Gbx�"�B��wM�IOz����7��BuU_?��<��c�{j^= ��Gq�|����F4���up�G�2�]*��1O��}�͎]4��H��l�o�Z��O��׾����PO�ۇH�
���?	Ģ����C�Y�\@����V�ϻ9t��DmV��6!�拟�[�3󄃮��Ǻ��%�H,�rE+�gZB����J\\)���%��a���S����oW(+Y�&��hM[�P?�y���-r��䥳���g��	�f��'��C�K��`�z},>����1���P	@��e�A_��K�Z�բU�^)i]<�7�Ў�Y�
I�c(��@�'pcR"Rx���{�@ɐA��.���-��*�Y��j��a�N�~�m�c�JZs����.�Y�Gu�� )]J\�tlNp�iY�
�#v"M��'�J(�$�Yn��Yu�4�\��+7����1���7T�@G��u��LGT�l��-D�$-������(��s�g?v	��ǭv �1Ąo��I�e��۝��6�5��[�9T�̬�&
�"�Z�f�=K̈́?A�!g���tÐ�mNu�S7����{�Ͷ�yI�v���_�T��w�82�U���Q'�~��)0�X#⩋��b��)i�V�8�M�;"�`Y�D�+�5���k�o�H�+�c�N�82���5{ i/�Rg�)�څ���Q@�Ne�!!4ݬo<��ߒ�����.�@ޛ��K���7:G4�B������t��V3����+�j�`�8�׌l/���"��ϲ�[T8��>"��=}%����	9��,�H��h�{�qU~����RC7v.���d�F�[����Q��Z"2�%��^Po�-�,,�>�-3��i��Fz��7s�m�Z�P�3�?�	f��	˙Y#
�3ao�I�TpD
��;_���0�6��=8RA�'�=2���ݚë*��a��[�����U���S}�8/�D�mM��0ȩR������aG���e>miL�>��X�A�f�|b�BK���h:Сe�`����#d�X�h�`t"���m��MG5NH���=�y��������aRd�u����+�s�k��#�$���FY'��H%�J�8b&������)��.դ���R�=|�0�q���-���*\=;����m~1���f!�_ܧ��Я1���g�UєU\b�&b���Խ�g���a��b���=��������Z^���#InH����fz�r�c�^	��_���c�I����g$;nT�Q�u�t�bp�{H��./��t�DXU#����{�<�FU4���j/�.36X���Ev����fh��_�1�#�c=�7���挌�uLJ�*��F܄5����s�.k½ϱ���K���`���7��8�Z��U4NX��W[#{8��f��ކ۱U�A��H���#���"S�n�����]-h��J$�n��۬9H��:6!�ay �`��FT���$��4�2��l�#��٪�'����hU�,/x�X��/�
�j@����M�v#h\�h�_ˊɽ�;�vO��U�Wu�e6��:���j���c#�!�T �*� ����1ۑ;����r��>>.���No���J��	9%$=n_��n�vǄ�B�O6}�{�� ��s��J���"r+{%�?�B��Z*�%T�y.��[�xUht�J-v�q0�P���?
�za�)���lK�:|[r:�:������)�>�RM��77>@�<W�pxCzR��o��Y bA�UB���^+�-��aS�k��
�-e�����ڏ~X��V.������R|��0��W�f�6\%��{���ռ�`7 ��\�p+��(*w=�6 7��c]V8[E�k�'�yn����79P��J�Y�B�+H��ğ���omZ��G�5�pC�L|A`�~���)����`�GP�:"����+&���p�6}x���}�' �&��9iN�t=�ۓ���+&��!�H5���Pz��H��!����k��<����i=��y��n�L����P�!.�m�{�Zk[DN�*�����tUm�� �K䡀T���O�;�^0*��������I���� �I?�/���4e�N)U�e]D��,g��x3U	0����7��<ؖ�	�Hf�#���`��M��o(�o!��	����%n%E�g�i�>me9$�T�` �U���l��)�jZ�ʍ�yJ4}���z�M,��>i�A>R�Z][Ü;	Bф�!�3lN�r�KE�M��,po+��'J�O�3����3łH8W7I�aV�衢q[1D	���k��.�=t������S��_�S��^��)g��'㜷 O�`)�C�j0�+��6o��|p����f.r�=�H ڳ�0�8ʥ2�PX�2�v��H���Q��9:�����b���G�W�q��X�o\u�<���J�*&���XG����G��fZmF�êe�@Ϡz�G�|^g�3n��B �bVvf,�I,��}<�|W�gn  �����ld/L8�&˸w�K����
r	���c���g��?o9#Iv�i�0$@&���Y�����T�s^f/94�R�hV��G���X�i�a��_[gfu�!z�x�r�!X�+A뾢Y�4`R&��;ZX3�S�,Y^�J�ŶSk����Ӳ7(.H)yl�8Z��23�ehC7q7-��6�o4�"9�1�쮣m�:<`��M�L��m����#q��RՊ���j[c��k=4��_�Gn���e���w��Q��?J5�'	�#��aNp(���ց�˿�1�+\@nL�h�m�J݀$5�}��!�Y9@ѐ+�)s:wR���Z5�P���@�1�8 �K���Y�e�4�`��H��Ģ6�� ����ڮ#���V&SKE��N�q"LAO�숩L	;4���`��� s�81&��������M�:���"�Z'����{I�_�wb��Ô���c�� E��o݈�s�9�ۨ����]�����L�gA1�d�, wR��ʌ��˞żCo6d���
��X0t�������K��xW��%�7`<��26d���[�u�ɜ�2�u���D-	���z0�޸�l���\ʮY'=D��v���t�A��2�K�9f��J~M���X�_0d�23B��xp><�!�g���Po�"�S ���O���)L�X��o�����g����`7~�7ޒ�q���+�������uU����#�;�Z8zVQ�\��A�N�N�q�07�����?]����R�d�&�Q����I��E):Z�O�s7(&0*�,mփ�d�
I���aё5iݾ�8���k����������Һ�}�aRJ�.)CM�Rڰ�7=n&�<������-op���Pք�GB�rպf��@V��]��<�ه`A���Z�_���]��oN��n�}E��H���������������a9s�������<��fZ�T/��MC�L�`�yv��q-���s��е&��r��VF�쳆�n@�O��x�]^��[X�/3�l���
��a
�%��r$:�gTY�W��9��!�<6�/Cc��U7�-�T��k����8��UEs�5z�庿��y�)���Aw
����n6:t�B�D&q�Z~�Tu~�~G���qQ=u���=�.n~Ԯ��Uz����Ϣ���)S��_�͟~!6k.ſ��A���1����
AV����ܧ�xl���{��8�A�ߏm�l��/�X᠌
	�I՜�Q�:�$q�b�2t=��\��k6�l Iu"�k�a��V��ς�)c�Og`�A�"�Ñ�k�3Ò��"`U�O�� �wK���RO2Ym�0JThy�D�ce{M���vJ��-�^���@Zg�G�R�-�97�5��2��ie�#쎀 �
�u��vH`쐎).�W-���Ŷl��>���������x�<��WP��z����{֬�\����(#�G[�1���ϯ�a�JJU�%���I���Fw�cr�Ac^�2RA��U��g�b��-��#�(��pp:���x+�I�%�T��=zW}Uԍ�>X��x���)��#�E��U�G�g"U��x��������~�Ç�؝{r��^CY��R�*+
Ư��"-��&�w|�OS0#���f�2"����.��K�hۛ�^=��T�\?���T�ꅚ��ֱû9 ���� �?�<�pN�&����L���Ж��u���)5��'m!� �D��US�%TZ���A$x�����	��
 ����=퉆������A>��N�vk��$ا�[j{䮙b}<$	
��!!W^�������O��QAS��4;3�P<�M�!�?l"��ӿ�.=-���D�F�~�2���~;�
�ֵ��M��Ҳ��Ve҃MB��&�X�p�w��i����珟��x� �Vי������X�肮	G_h�mM�Aq$�k_	���r��ֵ4�jɜ%�����-W
?�rdG�
!e�N@������+�y���`3��d�u�U����q�ԡ�Y�a��L���{d��$t�D�:±n�&|yk�
�ϐ�4��n�Pl��i*����o�q W��(��"�J� � &�7�[���;QȐ�;�� <�o2�����mPK{�*�W�љ�'�E!{<q�躁$q~����p%,���n�`�@�����aA�o��d��l��!�8���B�����'[��9���7�h�#}���!C4�bT�}���=�a:Z��{�A[4U�.=�����5Ϗm���́����~A��77��+2 �G�y����z��`�Z��Tg���,�)F�"S�qߴ���{�|�c"�|�1|�W�������g�(RF�7�(�t2���A�5ݦ�Q�?ܢC�<�d�wf���2��[�a��7O^�t���8�V4���L�	b�����:���Y}���>i�wGXDze.�HX`�1zx'7���)p�dy9<������"�H��yŲ���J����ڧ�!��O�V��}�H@.jO$�i��~�&T7��s&ӯ��'OcQ�\�ҥ)9����vp��� :��q=�~���k;�V]��g��Yi^c�jH2���Z�U�j���rt�_��!m�Y��>����:k�;+�ƊK'Z�$���(y��ӈ��/1���?_N��(1s�{�g_=�9p��9��b^�S��%
R�S��p�q�+������5�5�J��e�m���5m��K��3#�d�uKT�!s5�kK?'$	,�~����q�*[���8��,�9��+�9{�����2������x�E-׽��U/�@�Ͷ��|�ut�8N_�N�_"�+�����h+��%u~>���7��An�`n�e�qo�$ڂB+h���cU�M-�?��Z�>��-XH�UQ�5~w|x�{�[5Ќƍ��iq�-U�>�̿�q�����zT�����?�cZ�A�@R��L��� v�3e^���mݜ��WM ��mOh�k����,�)�Z�
n������MH�3^�U<m�^yz�$���ñN�1���X�h��]�/(�(F[��pc-�IY�ga˰�T�w��tQ�d!�W}��_�=��p;�P���P��*_R;׷0J��|�N�^���m�����9�6��]W�<H��s��.��D���|2<���X�:Z����)�j�ʏ�t�&�Pے��up0�m��=G��&Ӆ�m�$䩵}���VnM����@/�0�O^�u��\�Q�m�g(��#?lE��_B����t�N���������F���+fɥ�093:c��)�Dm�/-9
��l���~��h��5)�Lj\�m��a���s:�����=~=Z����m���ȢF�
kU!���C��ow�,�Y#�;>+�&��7,��UA������^��9��Psr%��TG-6�ͣ�Ӻ_5��{���jL�w�hGW��nϋ^r#�1{����L�o{��(�����B�wƬ�c��ޗͶ��j�i,:|�Bn�UvӺ�����P��Y'8w�F��
Q=���%!���45p�'�M���"Cߝ�ղ	^�Ȝ+��|��/>7v�9�� ��<�w�˷�j�B�d`Q6��ꀼF����!������d�\*`�WD/�K�
'�����f��L�
�4ҝig���س�J���cih�d��

��5�$�Yq��'�����R���>V�5�[�!P�d�;�b�O��g�'z���.�jO�c�*.�$XG���7���2�5׿�m��?ZS ��~t��C�F"%`i`%��IԾ슪)���ymSأ����	 *R��E@\bK���urG��_�-�	�n�;�c!��A����������J+�-�2�J�S1�V*�%�o�
�<�u�I>#IsK*	3�Ó��*�ь��~-�/��K+���Iq�fcypŜn��u��]1��4�/ ����O����ݿ��`ҠK��CM&�[� {!hDDcx7�|�і�jJ��������,J>a6��A�2��,��������d��T��bXL�no�GS%�O���GL��N�EBC���ť�%\5@`5V��V���B2ZŃ=�`�O����	�LA\l�Q���M�:f�O�5���y{<͋��/�n�q�h��tx
U։�mW�>�Z����{�{�\T�5$��!��|��p�����.�6%V���Z��~CԄHO��j��ʄ�c[Cި�m�ʪʽE!:�`>�C�g��k�֮X�n:D��}���"'>z�����9b��C]�v�d�p���r�Ƹ�I�ܬ�C�����Q�����s�Ї�5K�*"�1�S� �%ǋZ|u��-�o�k�r~���ֆ�r P���'�4I��a�,D1�k���u7������������A<ȩ��xmY��o#�P`��)ޥM3	?4�4B�,:§��p�x>����R k?u���}o���ɪ\*�c�w�)aFd�_#"��bWx�m�e^!pf]uUϣ�5����nR%掃U��_���=�
�`�� �q;J��u�D :�Hƚ����

*��9`�y�	T�Th�Z�H�5�+�:IfP[(M�Nsq��^Z�Q%��$��e%��܂�[�(��<[gsژ�mB��ׂ�:x^(@���F�9���la�]�ì�1�y����`f��b��ؑu����3�IY�5<���e�#�Nһ���'N6x�NH���G�	���/9! .>��Ċ�kDRZ�7�݀`�S�����#4���PU.����s�ӞZ,��9	#��I�'�ܕsk�ޒ(�����:n�k��`_���n� -�Jo�B��n>7H!�j�����6�*]}ht-�=�έ���D�K��t�0݄�"��}���*�N�	������Ɓ�7I�������JQ���!C�R��b�?D�ǒ'jy')�QnSLa�'��k4��R/?��D�\IS�{Ƽǌ�=�_�����?;��������~�?w	)��gx����v�ʞm��<�f����e�#�m༇�<���3w�~;/� �^�(z���`��}\]`z�b��8�Ʋϻ���^�ƾ+ͰM����^E�=!b'����`�(��VRZ�-:0ߓ�e�lT�'y�x�E#�o'����NR劀�!�*����3�e��DN_øߣ��|�f�|�A��h��	k"��q"r��=�6�,��S{�I�g_`���~CB��f�����6Ay ]VX�<��篏�2ğ���� �h�ϑ?N2�Q�n���34^���.'����L!���j����G
,~���J����qCT�����!�W�E���fۉu!���<�瞒;�t[���t��t�-6[EC��>m/�6��������>N�սN��m��^�2�[��O�7��E���p@�Z{�Tʮ�V�p��ŋE'�P:���D�P_�AA�j|�q��,8����{Q�}���t?�jF��J6�I�]a�F2L���Mڎ\TJ��X8c�s2���<�7��q�qz<��{1u�/&璺4E�P�s�A�',<C�� ��g 7��97�[q��J������Y�P�������!���*�|�!�0G^�����a�0����n�HB8����bb�:Z����-�T�`���Ë���JE�
E�n�h�b� �4M	f����JQ{'��JP*'��oə��B������;=��K��?+�7Af�� �s�p�|��+�Y�f��+�	?|Pq奥��jR&%�;`u���oK��(%�n�K�����F�A�*�|s���l�'^k)A: $6�H���-��_Y����ENRTo� K�E?�F�+$DX�4#Ǿ?����}'u�خ>�A ������w�j��,h�˶۬�3�Af�F@�Ռ|�?�GYJ��Nv�+�~����*A����!Ρr�5�ǫ7P��Ư�F��>NR��$\�v�o�X5O���VH�{�f2=&�qo�,1յпH�i��z�br`_���Rh2QlE7���ĐQ�R2� �|e{Y��ƊTSݰ��o�i����.Dr�+���������L��*'��'�d��\�ݪv�J��� �q^-��j�QI5:�팧���CY��7H��)Cq4j�_~�  e��C�`~͵��:BsVGL��Nn� �;������C2���V���`�i�ۘT��]�����d?���y���xT�l	�;3ch�����F�2�) T?3���a����nfS^);���	Jjh�Gm$Ę�fe;��5�
O���I{�E}[�)+Oڳ]��s�z��a	fv���CT��P̨8���ZU�T�|+=�Pq�!�J��;s[�v��0G��t^:�@��!�"Is�"=�!SS-�%��F�$ˎ����M���?C����q-���I�K��ԩ�jd�o��H��34��m��x��xi�78�׏��W��2�܉:��?�EI�ʣ��-;�^�P�py�b?Mʢ2�_6 ,[Iݖ��̹�7�ʓmaJ5��>�SiV��}ܭ{'<�B�e_%�#�C�8�U�Q�t�Y9"K��/��}구�e�?)���VӀ�pS�yx���,o";����$����!�;G���%��s����#2�=�b�`Z#�v3�=�A�ZM�51%g»M�f(�H=�@�}B�a���e�H�Ir<6[�Bv��q�[�X�����9�������.���t��"/�v�4����,�;���"E&T��B{������Ge����7��N����ę�_Њ��<�7�<cV�?&^B�7_�UK$�W+���+�ś�W8j�$��L ����W�;L����x�zd�aJ?���9��ˢZ����z���:�y�XlxVHYEB    1de9     850������j|�����8�EG��evd.ˎL�D7x;8�̓H(��Y�w����rw�A���(���Y�u���j;_�X���{7L��� �P�S���G��ap@t�'�[ӎl��P`:��W����,B�=4�u	OټkL�9�_2�~��z�����q��JC3j��x��ܩn��_�h��c����Ŝ�n���MO�+6`����י؅���h�}�A����� 3wcS�R%U�w����0�@���^�v����ߨ}3c��&O^ՙ��X��NxI�C�̣ O9��S0U��1*�Q�f�+>$��gA#�
qu�N�$|E�N�p��	Vf��l�+��a��G%�cp�}U;M����3�	���/�y�L=ɍ1�-�XA%t%R�^ӽ��p3w@�{}�����{�l\����_(����``w�:�+a�2T$�8ǼO��{�
�M�9w����?�*@�Ak�f<�I\S��"�$�����WP1�X&��[�v�bS���_�yļq%�0M�%�@YDUA4ŘRh�>A����[�|��S�O���\Ճ`�'���.����j�q�*��?�gx��(x�;�ˀ��t@ �z�$F�t�2�/��He�@�M� x^e���W%<i�������J� ��_*;�N\oT�{�(�V�Q�=�D0d�oָ�J�Z1kN	��^Y����5#���֮��}D�G���T!�s��A+@*�����h�Cr�S*�ّ���zCr'�=�H#��Y=������u��G9�o�)��wJ��R��`��d�$��kuW��� ����Yv��1$�o9����p�9$��W�*>�姓?ώ�� �硅�2�M����9E?&�B��dJ�Q+#��5U0��Ǹz/�72���=Z�ϕ�/�Z��^���<sB�!T��8ȟ�����r��j&��*y�!'+�9 ��U�w���[���?��g�%��[Nf�C����G�玦m���=T0}oF9�3�{�6��#�<�}v7ag&���H
�sW��A��R�4R��t�)�i%�n2d�-��Hr~���oo�Q0����ǥ�ZQ��iG~��I�� ��f>�c�I���N���C�#�i5�����Ș3U3q3� �	�g���`�]��8:��}�uȦ��I����e��� -{}49��̕*��rTo����5�8���,�����	��R�F�6�֟�%���`��-�M�x�^s���²��>��t�u�
ʋ �Z��~�Dj�����d*g �ç�r|2���nvWs�H�p�UN�i�xޡE�.���6�������p	(L�3�.%�A��M�'�9�7�Pi�J�o�m��-��QvBS.J�Z .̩�W�^�W���s���fpp1���;��bJt��t2n�Wj������xv��P�R��ڗ���s���?
Gפ�ך&�� O�DIL&8�^w��{��k�������+E��I�-ܬ�M�t:0����UB��=���)˵5+,Ɖ#ic0�h�"��Y_'R1�E��|�­B]^F���M6��Q�I���B�ū�&}���]��clx��W���W5�*���H}KJ��a(M�x#E����Qpt�����X��.݁j4aU��q���Wfh� �_l��,Ƣ)��X]Lh�����3�@�V$�!�VG��_Yq��~NfG+!�DI�ݖ�� �GqG~��`o�W��U+�<��%�_uJ1��LOL�p���?��7:�2��"���+��Zh�ْ^��J5o�������I_K� $�"Q�͊Ŕ���=������"�@�=#h1c����5��_����r�fۢ��V��ʛhݕQ�����܊@���g��Æ����JT=K4��Eݲ
՝	Imk���u�#�$��9������F�?�(RvW4t�"CwB	-�v�;�\���m�u�������ʗ)6�"����~�~�	i�'���d����ӽ��X�"5�c����LG/�iW�)���N��%���~��*����|�RK��&Fw�tW͟A:4�p�[��j"�z�f`�&ldv<_ p�