XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��+�e�P�"��T%>}�R���=�'^rF�z�i�:�����DJ2�@�ҥ��:��z�CY���ExBpC4�3��8��xm$V��P�蔠�Z����i*�����/�EJ�"�,34m�3���?@�_
�����4�;�9��t4�p�ju�-���<(wu%N3|��/��ch�X��S�o2J�v�a�̜,}����X��,�j��t�o���#'; 
���|�qD0�E�t��-���%	�V� ��'D,��34��bagλoC��\��y�F;�i����^�^�̤!H^�$�k'�Z���d�3�dgz>�v��	c�_�4<h���q欄)�6R�͟A�C%�R{���I�q�|�]�xd���}��n��������rM�ڥ,8�5 ˰�.5]+�f(�����f��#�T�[��kȍ6Rg�-�^|(I�Dd'Ʒ��뜃��$��k�Ѷ�h��{+r=JmBI���Z��|;�4�P���!9팡�9��S�hW��+�M���
jb��ʩV4)�e���ae�mбT�C�h:��ŧ���R�C]�kP������P/N�Y씬6�&�i����_���a2�e�Б����
��I�����^�X�}HqQO[���y 7s�b��(��|Y5t�����N4Ѷr�[�a0ll/y�������3�����E��g28����|9<�J���j����f�u����0�/yFu ��⽚���n�{O�D2���ri7�EzV�.�XlxVHYEB     8b8     260v�r�N�rY�lz�q�a�+A	��Q$yfHI���<���Ju�ݧ_����:�Q�N4���ަ���ʃ�j)��6��S�[g[����؅�8a�fƠ�&���ڤ��2?M�x)�#DE0����i����_��L5�|��܍ףh�w.^�����Vڥ/n,Ǖ	��',��-��샚���ʝ{��o����X>/�H[GZk�G�̄���ԍ��2�v04t���w�U��ڇgIS�f :�wEs�^q����?���*�X�t����������ů�躠v�맀Z����
��f�Tp{�]���[��L��66νx �:��%��z���.��;iA�$�9��,��z����w�����>ɑ#f���_Z�����x�/N��� 7�/�P���>`����}q�!���<g^�5�<7Va�|XG�g%�����W��l'�ڶ��I�N�E�$Vνܪ􏄯���pE!��t[�"�����	�����4�����L5�/M�/>�{�K����]���A4�-�91�x���{ �B{�b����/�R�lD�Ħ��M-F�u0����˭��t�Scbh�8� �-V�҃