XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���p�Miʵƛ���1)�EM��a�Y�H�䪖wbX�d۫Лc���tlGcQ^�Xq4`F��ݜ�û�X��CY���<�y�^5��� ��*"��yz����LZZ'��r�:Q�����'gҮ�S>ѳ�[��\�kGuɔb^8b9��_(��k
J�RCǃ��/�;��\�*�ם�'%�����޸*�6]B��Tr;;_��@U8$���l�d���3�F|��,��C�^�xL��/t�_Q��sm��h�\Xl�����q઻F:I�/b������߭+m�DX�w�=��BtXF�,�8���x&�E���J�0�i^ٖG�K�/���+NѾ��ƺ�
�w�u�[Y��Q��F�!��2u��K��Q��[�����r;��&�!�5���6|NG3�P��%����[�6��8n�d2vL�{[�G
[dk]X���)�ji�-|9�,�Uj7���xVc�A\�]��i0{�v�TS���!L�d�`�w ֝M�I+�ݪ��X���hZ��<oJz�o�?�VP�o�<�8c-������_�r/%�9��]_�[��}�5�+����ͱ��Gʱ�=��������B("Ζ# TBf����򑜑>z�i�Lx�(&1�*�s��-��UF4QN
��@�0[�;�I�.�������|�]�?�u��܇i��k/!�:���3A�p��_~H��QWH�*ǥ	e�`̅e,�4��P�� '��.敕����m�˸S ��h����%��O�:XlxVHYEB    2d65     c60g��/���C�}��QH�zE��L8�^{�,�nOK��3/.��e>�YJ*`�J��z݇�2���%�`l'q)�?�׭�GN�7	������ e����@m�R�9����l
�*>Q����xsA��3gN����/7q�O��j�<��5��W�L&c�r��TP.ĭ&�	�?��]�\|�EoeK��*�o���T*+c�dz(�����M�i�E�u7�SQ�H/�5'+K)9?k�,��h&Q�9��E)?R:ͼߘ�8��6�����GȧZ*��j��B�W<=�R�Ӛk�t�Y>u��l�c�����T"�dz�ZaI�9�-�Ss��������m�nZ�+#��]͛��8�Z�B��O$�.ya@�ǡx SL.��Pɹ  	e�ctR��_���kbH�<�R��O+#��%���/�����~���N!)�H4�hpgʭ�W���Ό7xdd'�I''�KL�-1�A�3?@]+�'M+�Oy� ��=e��|<«���_�mg��jT�.����<�����7� �"��&�`fM?K4?��������"^�]��ۂ:)���ٜ��]m��MJq/���X��s�O'�XI����(�.��ъ�`mjХ����H�2I� �<�~7UḪ�:�y��D��~1)�+0;&9¢&JY�Ǜ� �|����m�gO. ���D����9�QQ]�z�lz�����%�.��(�-�L�>2Ito��3R��E�J�!���^��QRx����;���7�I��/R(�4VIi��}��V!Y\�!:jB^F�G�~ ���Y��Ys���ԙ��}�
EM�b�[��1�����)C-��]^ɇc��ϰY���q�k�|������ۄ�,�B���~��k�Ȥ�i�8/�S�q�S'h/�A�g�o/ic��	�V:UD�!T�M�p��0fi�i��VZ�-G�ĕ/��j����$̦�w����f�em�:�^n�r��o7�\�mf5E�Y;�xQ��=pr$u���q�e�0,n@���ߝ"�3�X�(��" ��px�G��}���K�'�6K����]|�KBo���\ɓ��_LD�L����Z����:��{�DZF1 �Z��+:��%Tץ���\�����:����;dHe�t�<�QS-�cG�1������__CV��
��u�u�APbNy�_�[�cIb��E�Gr� ����W@�km�t$�?��UV@��޵`�y$ y��wG���2��]�}����T­D�r#�/�5Ӄ�5���n��E�|�l��u��4	���mP�q�T���[�/���W�;�pȔ�O��M�9�
_p������(��zL��4�?�5�u�̂����'�`��@"�D6���nW��6Џ*�������K��jE�/��7��\���,x����#܎)0N��6rM.�x68��,-�k-��o��-��&�mʉ	�1Ԭ7��O-��s�n��5wv.��Rٿ 8�6�S�H�*�o��jS"�3�\�2Biy��j����'�� `x�B����i��!�P�SӒ:A����Z��W:k{��o��=�
T��E�1���,~��i����zẊ��_�Ф��ޭ.g���p�
��i����ʂt�=9�Q"0I�U��K2g�Y�(@য়�J�����$W���k��4�g?8�Zs�h��MR#�ԧfo��z���%��a5U� �*�Je��� �֎E ogt����ݢ=��J��?�D*���C5:�
��R�iL=I��I^��kPzǙ= ��j��C"�����˶�����k�v&��C{����@$���FG�eBT}3
�=C��p�YQ �d��(��'0U'�"�[��U���wb����w�ܻ�Ќ����&��ϼ�.�vsD���~gMAf��|-��ĝ�*��9D����zɕ�&����'U	�a^�1�2 ��X���?�Ѹ7�'f���<�&���H�F�������[B��	�Rf���OŸ�'f�P�i"�kx_ji�_"ʦ/�7����~�>��=��$�6���.���*�̚��>c��Mw�L]���eP�W�[%G�A�i��� �y�Ț�j��n"5���n�>.<wd��q�h>�F�.���Q��d�H��r��"9�Fv��v�ZV����:P2@6����pO�+#�X�H�8�^Dx񚺦H7,��>����ꭴ�R���u�����89�F'�Y~ӷȠs9�	6��
?�� \�?�!���!@=R$E�s��d�����mi�W2�z
!�Ժ�z�aᣩ���g���^"l>#U��P"yGw��@IJt��x9���|�����m)v�E��\�����9=~W�A0�=5J K��-�1��[����2������S�e2�Ϻz�)	�4�GA	A��� ��&�Ԯ�o���N?�
Ճ:�<6F��^��q�Jj�i3�����#�Q��yl�PԞ�y:� �p9Yb����LK�ꏹ�΂(z�1.���B��w5�m��!~L9���?���=���I��,�����^x�#�����R�<����L�5	�o�����{H����p�����6Հ��B:�@1:��Aʃ���p�}��,��ܧ_z��4�i�wp�@:�\LSӑ���wu�JZ~�)�my7����c���C����d�q��*��P�t"�K���2���#�(?G��i���L9�.�=��SS2����i�#w��0��!��s�[��E(��_�̴�z�l�F�9r�������<���/?�;��w��^D�/�7�k��}���c�A&�nT� �.�yg�>�zQ�<I�)�H��C�0Ȁ���~'2�Za��Ň��J�Sw����>ƣ?o �e1�9��׺�b}M���m��=i�X�$�&�W֦燰����	�����5�ĠD�G�n�_�Y��%��n�{���Ak�5�ɢ2I�#[r\?�YI�  ڛ���=����y!��"T�p���ֽ�aTVg�˯j"M&7h-U�?T�26%_m���:�����I�$��P��KB���_��T愓���e>p�F6���[��@�Ƅ|w�B�\�Ķ�W�� �,���s�<�=���L���f�