XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���yָ�����1%��+�~g@\�{�+%,4DAD&�m	J�c,-�
1��K
�Bsws��� �<���z���m�2J$;�P��é���Իu
B?�,���P�٦@�R����M�ܮ[u;O����&��@�N`��}���DGu.<5>!2�1˸mB�v��jUk=<��D��JrȻ�E���2]S~��-�>�cZ��7g,`Z~�`%���v����z���V2�����Ch����r�R)�b�}Zm�c�k�t|S�h`߱ ������&��Um�n�\�������Oj�xΝUJT�0��]�}��$����k�Q&l;�(v�㴧v�sY6�c��&�P;FNx��}�O�H�_�v	C�K%��',�<���5���U���w���r|�>����`^����y��>��>]���)L�o�'Ƿ�V�yn	;��*wβ]"
�'����$��Ҩ��ɱ���U������zZ�f"�9nK��5Db5l�� ��~-�������9���mqdp���VOo�S���r�c�[�j6�Uy8�-W�[Ԉ�&�>_(���a�q��J4t�1f�L�/NuW����i�5Ȼ�}����Q�(��	���yB1q?�R?3p��P�&������I7EO�J�ƚn?�Y^1�����Z�;��nI#X�AQ �>���WX�]Η����,�j4�Z&�
�7��\���29.��:Ғ#�;�ʏ`;�6��v�A�}���k蠃>XlxVHYEB     590     1f0Ѽ),��J��E��!�g�J��nuվƝ�ו���Ĕ��v'~\'Ec�n�c���n��_���j{n�1����կ��)��]`�ح0���맅�}��1n`@���� Zq��Ɓ��`??�LCH�S���_��k��.;E<���a��<�iO-"�{��C�\H,>�!B�!�{�㈈�4	�>�7#	��'���C����Z0**{��j����c���|�;�2�:(���KS|���^x����P䎉t<k�F�v��Q�M����@d��{��8ԋ��VG{��ꋈ�t(B=4WqgOH�@��x�v��i�H�
�eqD)�g���+����崤q�UU��e�'pQ��E8���_A�A��c[�Aa"�;SZ;���uEp��oǫ�M�z�L�o��1����ޓkNIc6�Ҵ:M�P){�;�Tl��_�M\�6m���R��T���h�Bn��%\{D�_���wp̭Lͨ�M%