XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��r�}B���$�Őlۀ�X-&	�6��(?y53`�>�{��ޜ���\M�
T+�C�c��K��O��"C��p��D�����b*�ȓ"���5��5�#���j��@7�Q�e�h<�v�?F�=?�j���u�ns���p��2Gz@� �n�X�@b�aoV,���/�b`r�E��m9ْS�*=Qmx0;x;ǖ~m�"Y�5�q�sp����|���/$?�-3((u��Ԝ���G��[֜AOu>��VT����b��������;����\�"4�ofK>�C�x�%��|��Kjԭ6�6?2�2��[�����J���|�"�<��|G-�b���& ��^
\�m`O,�����<1����iポ#0��e_���+�=�,h}�߈]����^Raz" ���t�Kć��	t�k��+�({��I|���$�����^���M�H#'�
T��е�>�e���hr�i�t�����&�<ꦛ=�+�3�U׼2o҉�|�#'牬e��=�Pv!�q' �%�H�����x��T'�¤
����Tp�Κi�h���C�`|��)���!��{8a"�����ݖ����I�����d���O�����%$���r��l<!�\��\+�A�%�B�?R��>kvq_�� �ʹ|�B�H�����5p���Oe�Zt���z��,�>}��D�7��֑�a��yh��BL�g7Z?����̧�˛q���Yt%�PqW"^���{x4*�����U�8l�XlxVHYEB    1560     8b0��N�t7b;�US옫Pl	���LV\�����(p��tP��1M�}ǷS�f��̏YU�X���	|j���ۧ���q`oP׵U�!���+���c,U�J��4
aS�a�=�ZL�����8*K O�)˝�;jP$���U5;���[.���>uU`��x���iq&"(\_��4@�'�ً�j���Kb	}�T��v_��J��[oN��s����x�v�������l��}ù ?�^a���Vgf��Զz�ɳ�v��	��M��J�3��c�mN��ÜD͸n��?UWǗ�\�N�������,B���x� G���Z�3�Y�XR\ܠr܅&�̅f�ήM�`����CQ)��)�!0V����c��e�Zi֣���'͖i�} Q�L��V^do�"��@�LHl6eg/��2D�&ኵ"{=�WtM���/z�1�l �G�U�tH�@�Hw	Ҝ7��=o��6��\�+��p�DWݒa�&��f׻3H����M{��b��&A&��
g�GS� ���eyHe�X�Nq�ʼJ�VLa�.%�@�H��S�	!�pΑ*[/�0�D�^̔e����.��@��jos|A�E�->��o�P��<Q�w����`n��TOd�5KXk_>��xw{.�������#?D�i�p�5��4]ߥ�E!�xьۚS7�)�^����@(���� ����[E0	�U[u2l�~�t�otS�����cy֟� Y �bʜ��Y�����d%�O!��ʱ�zHHn,��8��r<��"�%-#��q��r��`�a����A6n�n�tӜ��c�`
�on���"0N��]к2�vޠ��4�ǐ.�T�����%��X�M*ܶD� ���V�N�������YǙ��h4�B=�c��aȼJh��0����P���ee����3v�<N��}֒y���[Cs3�~g��샐����.����Ze��pT-}}����iO ܉��y`?�`�p���G�.Db�'+|���M�L�ݔ���R�5~���Rd0����zp7NU��6�uN
��$Ftf�<`I6���>����@�
���yi��x'�ƖX��!��J<�1;��ĿhXd���Q�%�p\�`"E���o.���D+"�5��
uu�g�Y!�ԖW�֧���7]r�?�P��1��V8�0]$�������ύ��T��������տy�#��Υ�3�~[�Lk�˽T�<��O�/�� �	y��֙ٛ`~�FI�8��۲�Ò���L���G��O�o̂����*�X�"�_]{t`Y|'V�ƭP���v6K9n{sxh9�*��tQ�p&O��$L���/��D]��ϕ���N��=_(�E�u�W�������	��4��Q��e[Fh~�KNs,d
̎����{�U��	��;)�/�s|�[W�ij� �K��j3�i�"�q�����IXF��ٻ��z�5��P��!:�������V�F���z�
X0����:�㞥����U�*wm���8�xQ�x�Z#e�'&�d¨�7�۷���=�b8I���ѿ�AD�a�PzZ�V�N�9�Y�C�����<�Ѿ4Wρ���
�ŜK��T:V�
�j� �2aZ������뭴>���
X�"��2��`1�sZ=�����'c��4K�ب�3m�@"+��Bx��'K��+X���5�h�g��$LŝO�r�Ռ-�8k
�Q��� ă�&V�:�0�+Ҹ �<"�A |	��߳Bf���n�x�n@�{R4D-�P��&��g�m)5�=kbT+�ܸi���q��.�|���̟�;"7Ce�C�R���˜�'�E�U�0�A������	�P#��˱�����9��
d�*��s��P{Cg��V�]�q5�Lկ���Ew-e���
>Į��<8O�1�s�a��g�6���w�l��KÙƽl���/����<�/lS�#�{8^H���?�ٓf�6�+��0(!�$��>�f1D�W�C�+]YDmJig���Mm�v�U[��ww3�0�gA���bġ���"��f�9�.���v�]"��Lh7�o$>2yF!�A+��"7t��-�6<��]�y G<�~��3f��L�:f	��w [�l!i��L+�)� y�1�,�c�J����9Zp�<�-$6��Õ��3����W���C|�'��s$��)S[��L�WKuV/e��`r2��5
��[;	Y����	�