XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��&���S�@}7� ��=����o������bWi������ )KAm��I�L�H�kWftSB0�;�:���KI��R��[O���@c/=C�<fx��R�7,�r��Yl,��y܂�!wk�1 $&��+�xY9��&�<�A���/]��lt@ e�@7�-���:��l�h���MF��\��8�d-4��M��&<�M۸��R�Ǵ���>��m)��̑��܆G��X4��L��M`̤��us݆���d�E�%�?>k2�Cb�呗��C��/$9�E����v�,��;X���D�C���wۄ�4��6(Ͷk��:y��P�f��������`��tʋH�ޏ*�ﵙx�V����(��P�&?�a�^L�y�Z���뀦�0p���o�Oqz-�B�^ܙ�RT!��#�X��!Ђ�v[�N۵ݐ�7^�{���q��O�0uZ=�u�S@*�n������^v�Z	)�G� Qe8=A�"HX�/�y�~����(ݺ`/w��}bn�v��b�Ƿ����Y��kR㘂�XK�؜u�V�H<><<D?N-R1X�'l��hiZ��0� ��U�<�"a�0��R��9IΙQ�!���6��Fj�<Qݩ��KḂ*�����dzF�ﾯ��6I<��p���'�}����z�Z�����V/���=�0���#����hm�/�\�c���o�p0�і1���]�8���k G�&��z?%$����(����+ºg_J�ᆔ�@�XlxVHYEB    fa00    26d0��Z�����6c��+��A}A�&�#��1��&I|��%��{�f��M'�V0��آϨI����!h�gAa��5�Vc���`9�{Y����d���.y��}j��ɩ��G�����$)�����!~/�uxF���2ny܄��^MG��B�<�(��&�U+����#�Y����!�����wx,�ك�\��zI���D�lr� n�w.��S�m�A����_��;g��Ɠ�X*Ҙ�QՖ���%J;���ş�Gi�$2ҕ<�	(mxN�[���8�ĺ�Y�-&��:�F��%B��u4�͟Ь/�KKH����	Jkn��!R�(Vƨ��q�m���{d�K�G�)��Ҝ�Ӡ�Y��~��"��C{�X��F�> 4�����˱�~���r�]�MaS�b/�'��O7�X� ~���:'F��M�V`����-o�5�\�WI�.�:�G(.ol�G@���S����1"@m��eZ��
藵f��-������%��-ܨ
���od����{���QDz��	}Ss)R"*�K�N�`N���T��L��kQ��ưN�s��ky���;:�`V�}E�	����j7�jl/��a� -���t4�U��~�4i���i8�I��)yk�_l��G��lM����)ń����	W#Ƌ�%�!�F-b�5���k�0I����r=�&�j~�I��%q>��n=��i�^���#~u��q%&���2`�t$�9�@�9����HO�~���������E9P��m�[��~�m��:M�="���~�V��^><7j庂3�K#[�0z�b`���7�}E7����%����=^cH0FCVdb��e�[L8h�H�Y[C�~����<�B�}�I����ȴ�-A�r���a��凿N��M��FXKRv7�MM9����4���.��l(��(9a�>Ir���]czsQ�K%�K��Í�o�f����B��_�U_�J���_���&Vd� ��A�@�+9������a�zṆ�ᕲ-Β����E�|ٝ�B�K�t�⊘�T��U�����	�}A�l����x�m	xE**�aZ1��]�y!�y�n}�'��ay	����a�0w���m�6LYV#:�GQ�E�:Gxg�[����v�r�>���*�x>�Ăm�uߎ��lF���I8ګD�(�9'�C�tx9�An]	�57)���Ӟh �IN�nO*��t�OƐ��;q���T�>tC_��P�<5=v��u��)�����3�`}'D�����A��1Wdz��"ݑ�z,�o���a�l\�E~�J�[��y��_7�,�E��5�4j�
�9���b��M7��ݵdg C8���Ϸ$�`<�e�g�)�xdy7�D�'_Y�1��.�τ~>���J�29�%�	�.�}^�u�mEE�(�:Gb��,U�X2P$���[��?��1��[O/K��kf���Z�ְi����=veK&%uZ���-㕶��#��ص�x��]�����0��g����e������|�7��гDryE$�eq����S�T*i�u�&;��_���`����O��!��l��\� ��� =���ҡ�X��i�a4i*��t�d��^.W�����(�T�>����������.Ԡ40ln{��uo)�������s6m`hUB3�׶�gɥ��+�ߞ��W�K�O�@�H$������KqSB�䢙
ap�4$��.��p��a�C��:"�#?/w��hnê|%�"�(`(R*o��;�����|{�=������;�u,A��Ƚ���3d�|o�� #s��S�ʉ���IR8_](XV��f����-�2��	�j�@?�3�@�O�}�/Or*��17+��_3���$Q�[,�X�f��;H����~W]`	P�1�
��l�(p���ڐ�r��TU�*�e� w܍Of�5-.�r���K�����	�W�ՈpF����,#5��.�sC��y�Rܡ����[~�G�i�������n+��r����ts�f��հ����Ӱ�Y�S�aT��YalN^RT`���'�i�~��K�(�W�٪&6�PK��A�Fa��f���Ե�R����P�
y-.ђ��b��Ϲ"ǁ��і�e������?�^�E�U�a��eg-��PU\ﶺ=�m@K���j���-]Q�$��l��~��q�@|��o<>K�����R�3S�#Ղ�X� C(.���V��~����?(
���(Xi�QҦx���{���ਗ਼l��''9�� ,>,�1�ߜ���S�:�Bh� ~��}���t��~3&�AT!��`-���x�L�Y�vLhت���1�L8����G�z�?�vu����� ��
-,�<v���W��x4{6��^x�Rm��V�7v��(h}�����q2��/�%ka+2F@�~X�Y��,Ş8'��r ��dV`e���˚� �bK�ʠR�S�ͯ�,��r�A��@�e�꓾[����`l�YHr: �y�,�6oGD�d1�k����[$����`_��u���,���Q�Y!g�l\U�AB���EĘ!���v�X�b8bF����vCh��,�����z�����	�F�'�!H�(���8-�QYqJ�����( �l�ճ�������4���>��!+)D��o77/�4A$t�2�-I6W@֗g��<��M5?�wP4��q��N�>p�V�%���u�����O"�"t�֯1@b~
M�1b�sn�LFt���KQ[���?ښ���nH���xt~��@��}����Z0ت���g���-'ד�_D�R�__MNO��uIT�Lr�[N�mr.�ڼT��Q�5{z_u!�/�Ӯ���� @������g� �+Ɲ}>�Q���$�R0�^0���3����	J��݇��&? �Z̠�T�G�-/t���,�t�g�*}p�;�w�#������+qr��pcb��U�~}�?�cV�g�}� D�<�r�ē&�B��ۛ�Ec�{^�O5��F?�0K��f�T�f�����=:��و���Y��XH�7[E�۟^��=�|1�*Ըm�K��,���&���t��ߐ<R�2J	�� 6 N��}��bg�|�D��Ó��oDaH��c�]��A�ޓ�v���$�e7ӟ�G���Ƃ]M���,Y�?�ꁋ&'`��X��Cz�*�@D`����W�zE8���9�h�/:߭����?j��=��W�pm�����+=�ڈg%PbΈ�3ʹ�N�Bg=4d`�
�!<�F����|/���f�dc���(����a���:�*8Tgq>�c�^�ϯ�E"��KXArjJ��2V��[lЅ^��k݁5,�%�R�$��LxayZ���dd[[H!\��uAºE���������n��:�b��:c�w2:��Ե��((����U����.V%۬���&Ƅ�PN�#dcX�F(܉����Q0�z����8��٢y�?�&��{�g5�c�Z9JkЃ�Y����Y�%��>5�4���{��R�P�<inN.,��*���UIGjN�ԭ�.����bu��y�P�I*"��l���z�g�p�\��0��Q�QR��C�!���9�_�ǜ�V��ɣ/Pޛ|{��P0��!
�Լȑ��.٦�U�a>"�����a<�M�^��ҹm`H�|�f�<�@e"�ۋ�N?|�S�c��؋�G��v�޶�\�έȱ7H���Dy��.pC�喿y��g�Ml��O��F�s?
���$�,1�a�H���j{H�H�����i���e���-Rk���f�5F:�sTm��Πp���zSjm$�����5�G�u���Q�xܠ5P��J��⿬����6`�Ӫ7���Ϋ��=�����?�������x�x�a��L^v��l��>j��%i��V���j?����$IS{���9 ��Jҗ��ݍv�I#��g��f�l:;��p��(^�E8jܐ۲��=w�(�a�^侗� C>Ġ.5�g�f|5�E�N�#,*�v=N�A�_�|��T��(낕���l�>#��q��ݽ^I�
Cu�WA���@�o�U^RQ@��D���J�&�8��Rߋ*�HR�Sb'��D{9����$J��;K��\����s2�U���ƢnH��9#���@���±y}���h�Ⱦ��M��i5�U��D����[S� T��l���v�8�w]��}m���`�B��Z�*0��{���LNH�<����P�+��.�A}���s�� ��Z��H��Q;��Eu�c��dD�D�a��i�$'��P.�h�TO� �G��eFyY�ٳP�&�#�8��PC]�f�#"�lC�3�2C��h/����BpL���\~يq����8q _�."ߘ����gE�RbR���eVk�3mܹ�p��F ��1)�N�䧉)a>��îG��Y��<�^���j�����?)Z4'�z��Β#��v�O4ht��Go)� ~�����$���1��t�|_�����8�Џ8���r��Y-8(��u����\��
yc��ɿ����C/ ub���lVk�594��[ӀC�)C�Z3������N�0wҗ���3�I�ʧtT;�c?���K�j��!_�Z�;)����'B� (�l�>kˌg�W�|.�P���K>3D�K�կ$m@OMꋡ\���T�*��7���5�����R\�h������ye�=q֊��1؈&�)Ǆ��������K�"/#�M�~y��Pڪ�=��#+�)Z��%޵j#��v,X�{��3�Ч��ftM���]Z�9�_Ji�(����A�%ɕ��_}'��������|�^�O#ʺ[W�� �Z�o�F6�����T��Yz�훑�Z��j*_�p)�EDfC.��aF�>W�ų|yM�{�5�.��&�wܪ3�p����=4 0����m�|�?]"���A��°��!�!$���-��&
u��h�%:&�Df���g�9�����ߦzQ���qeSË��D�-Es~�t��;���!p��/�u�aJԾ�Tn�)!e���p�~K�����O�eN��R�֘4&�aE�����'�ƁCp,rv4 b��r���m��U��N�z�{����̧b���;#��(�׍���|Q���������CD��vW�V���օ1�3����'��
n��m�PО���ґ�w'�m�m�i7[����sy媡�q<�j��m�5+�B���c,Z�2M��mـg]+��;�;j����شw?mF"��E(��Q��Iݾ<:Qʴ�V�Is�8�q���Y�ԃ�4y�(g��S������$�,�=�\��	��?*�t�7��ۢ�GF�f�?�/�a��n�uZn�/ʡ*�4�"�
��+�'1&� ���d��J�bA�/_��:S��6��1v|[6��k�۪2rE)�\������\����l�& Fc��g��(BMo�^
�,zZ��%�v�$����\�齕������E���_5�'����I�Mx���6
���O�EH�~!�8�uj�/w�q�j�˰�W�M/)'8���l4N�=: 2�J��;&V�X ��߆n��e�3}��x���d���z_���})�W%X�v���T*��y1|D���z�	˄0ja� i3��,�*���� �t#Lpi����֐_������:�&�����P�*����(Ƒ*A�M݉a�n��eIT�)/x���V���1J�N#�uYP�PDLS�q�E�u�IQ
�e�U����.� ��R���@N���Q�xS ��#zAaS�`ׅ^�E�\	��ϋ?�ڻR
o�9\��ǅ#P����}iEDԏ���}��؋�8�r�=�Ɛ도�z��Ey3��7kUz�t(�ͧҳ1V�!*�n���t�؂"k���,���Cm�����q&5���k
;"������0q�" ��> Z��j�+�tx��C�F����f{�0�����0Hƥ�2��N���yQ`,$���{��q���?�%`�'��IH�����H��b)Jj���p�ڗX��\� ]	ka��li���ˠF�Ä�o��!K�qs���z��*�@�0�[x�>�g��8����hy�N�;4�|kܮ
��a��1�:@ogU$��%��b��_���Q�xn�3c�������8WY��1��Fx��=�}ݯT�"��N�_H�N�=zד*˪����ҳǬ�勡s%��X�d��R�mn5�]�Q�^i�}pU�5e_��L�Z�hT��ܟ���D�l��^Pa��q�EFh���(09�|0O
o�\�u$ �,��6��b����޴�&6�9¶�FV�	W��4@\I�B��4��6���֬4���o1f�K[��*�Pb�z����7m3s?���m<�)��X���������ܨ�[��ג�6��+�-���@��7�������Ě���M��򁢶�~��C�ۊt��G�@m�1�c�l8�tn�Q�G������ȪH�@ �c�T����X����p�#a6�e��鵠'��<AqƂ�(B���@�{�%����І��ID$_:��d;ڜ�]�>�RaI����	�pv\����{ =�n*�י�d����?s���)<�ij�@����������� ��5�!�XN��Z�aˁ^�l�R�[��K;o��q�_fn/�(�|�����{�'SDtO��Wŀ��m��%�u����n@�ͣ(���KO�Uz>���2��)����^��I�F���N��:�y�`:u��tm�|�\�uw��cƣ�`T�
�k?���������B���yĹ	���W�[3<���	�{{$�[Q�4�������
?)����rŇL|�+������8j�y���z���^-�fU��b'�'|��a�dv��!ZZ$l�=e�
#��k�����H-YE�g������d+R@�0�� �d6`�8��LY��� ej=��7b�؅�*�����$u%c�t�Xgs%����,�Ë��{�z��҅	�Y#t9��ᰈe`�Η����(����3�ߦ<;�X}'�wT��Q����<��`K_[���P-A��SQ!n��ՋJg����^���-O�F1)��<�i����--	�^& ����Kb��
�m��{�����Z)+Ι%СͯG^��uu�n+_/[���g4�gWJʙP؝q}d��=��>��#5�@�i�@�$2%w�W�D���)
�H�JÆ$',�7�Y1��N5���3)��A�:��I��'�{�,���?�RwA�so��P�my� �99�T�p
�"G�%^��gr�e<$��H-�9�g��M��&�o�"1�^MB�I�����32��e��O�'S&7��.5)��q�:���S�d���pt2J���p��6Ʀ�]��q� �����J�T�g���z�^?�q���G��<	���-�2�1�(E��V��ʅ�/|)u�7��XH:T����.�yeƧ��ݕ�4��#�� ��%��p���N����1��o��b� �IG� ����&h&�!̱d��D���v�B?\qh�����	AY�������|��z;$�xH���J#��G��9��k��+����&!�}N�\�ɳ9a���*����yަ$�N�wLW_�t-��'Q� u9H��u��V93F�E��_`\�]���.�u#�	�h7�Ϩ[&Ǭ�;ЛG�*�(ߺ ���R�%w6;���u�X�Y}��K)α�uҬNJ~���}�k���ΤpiB�'3�Q�[�Izk�DY��n�H�7�d.�]��(גl>C�1A?r ������=�*7�7�
T�_W�H�\\�����"�D7�Tf�O�\�d�K�WQ�8<rt�H�j��؝�S�|��~W��w�q/N�B�]q�M �f�����_2h��0��A��}1MK�������b�c�]h�'}�t�;+h���ĠkX�z읣���+��)�0��5�����\<ӰRE�`��Ӟ�r�5N͓����Q�]�I}�%*�ص�lC�O���4�ܧ;�*�ᖒ�b�`i��f�пv[���Ij��QLqe��$g`��Np�/\�	��u��-Ki�^���B0�n_�O|�L��W�_7���޾3]�+���]�$퓬�؏rs���
�J�~��G���V�%�N���pBU�Ҁ�-%�T���O���D6�$��[#=���f���3�����N�`�
0h�'����p�	2���|i�w׊�y����}��7f5��CuG����ن�b��GU=�'��g!�Ğ-�6�k��/-��O�d��&2�!�h ���R��ѧJ�Ĭ���wX���O8|X�ۭzlRːYE�RZ�SbEsne
]%@8��2�7�W��;5n�������f�d��?������/Zvw�5%��\��s[������d��HZB���+�g�����X�O���?2H�~U���<7w���xzzS�ӌ����Yl��ښ�O�?J���t
G������e1�����bE��r�{R<�W�_z��S �U���l�YTJ���vC�k�%68�����g��Kw�]a
�4�b[�6���5�Tv;ld,��֗�(9L� �Wm{�&m!��WA.� G�f#r|D�B��:Ǜl�5ۺΪ��[W�C�1o�O�k�0G���s�fE��>C`�5�=���[�H���Ow�0�f��Z;��Tf�����Tl��}�q��yf9���=m�s�-�3�U9���(\��*>`�n�$�lO�F8o8f嶵x�r���6r�U�eE:�Zߐ�#��gA��L]qY�Gx+Y���D07��jec�1#����=:Û9~�p:�&KS4O�=�R�D���A\a?�Ox<C_����K�&��D����}l���C=ي�o��A�����6I�?�Qܡ^���g/��E�t�Ul�;H�CFeTD�8�7��T��N�TG�V?��Z�kF+_��NZ��`��ʙ'[��r ��Pq]?���`��-6@���Ruz`�$=�8%��,O�vb�������7wO"���\V���vX�O�7�h��70���ht���G��~�1�i�=��w�1��R}e��Q�@z�v~��B>�h�ۭ[��M�=�h�x�d�':��B>�w�&,�����A�vcHY��!�xm��+��$ƘY�,���#�t##�kSGJ��ƿ�[�x��]]�؞�b5v��ڑc���szߔ��kݨ]M���A�V�� T��9L�4Z�r�T���]�hs��/ɖ\��z�u5�����-��W�o������85�&;�0�~]�4i;����&�w���T]���P��V.�b����#���� n�{GD���a�Xi�*�f���'����B;�Or��	c�UIJ�^��4�-�Ăw��6��� <Sgl��崞�F�C"�.���b��6�[��[چ������>ޭ{#�2W������y`��3g�Fۭ������`�2î8��/no�y���{�H��:e�j���8���ɔ�=��(�O�G��s�$�]�A��=N�Z����?��@�TT�������"l�u����I!���z�OuM{'%��3�S�lL��E�����	��(x��F �'�!hӻ��N��z��.}�o�(�K�¶N�Sͣ_M5�ySA~�`�A����=�E-�����6}=؋�݃�	*ƾ	�XlxVHYEB    fa00    1050r����د���n�F�_��hNt �/��[��S�h����^�˸g�1�Aff�U� ��"Z�r��~U2���	Cmǌ�!1]6M�t�jB��S���I�[�h%r�?8��ڍ�����	�������B���Y梠}�Z6��h����ӟ�9��ٍ�V��q�eiD$g��T�[	��˸ĸf'�Y9�?�O��+�F�w���n���� x0`�?�R�L$a*�7����LT-Hpv�k��
>���MV�����4�G)�`}�
�s�e-D�a�ӕ�����gMksi��������]��!�n�]/'c�k{�Y��h#��	�8���T��*�P�L��Fw?g��tn?�(:o��'z���'�6�ӝt#�[veU?#<�A�=fR<((D��̦�I2�pM ��9X��uW$���'�>�4�h0�e��+�)�P�㔩e��
q]
�i/?�,eU���=θ�&|ٕ����U�����5`�0A3��쪹��Y�0�D�&6c.;��jJ������s�Iv<4��F��p�R5�\F;gT� %���BK�i�Pb�~lk�v/�K@} ��]�c��J��ҎNP{�N9���!���j���я�"���r?�yi��m�{x���"�.�\�W������(n�Wdg�(K��ʀš}l\�W���T��w�l���sG�1�H��}��� 6*e+���7�.����/����kn�.�A��ن�j9�y�@H�z���j�@=S;l
�e喂���y����l��	�6����RL��Q�r��@�kw����;��Q����59W7��Z��z3/S@S��R�ެ_���~���]�<\l	���hB3��-�M�;�V��7�#�f}r�
��B�BJP@�����_���d���o�̭kEĳ@F����J9�$�~�:�J��~����̩6V��j|ǘ�p;�	f�Y��n6�lVG7R�����I�Q��A�fZ$A�R�����{ы�˼S��x(�h_��$�\��gB@�x�=�,]0c=nz�@L^�О�s��c���bk+�sK�Fa�,����x=����9/�+mQ��EC�U��/��FcBi��l�V�`4��	s�܍V�X��?����r+7.mH���gN�e�!�a��.�&8�g��}�F-m��0ݫ�>�̌����%L���9@����˫�[�sś����{
%�����o���uf�1�&K7���� �T�~�X�A�� �n���C �FPT�
9Ρ�V�m����R�*����13��+a��_�m?��ߐr��F|��Ep��LƁ�	.Q�BĽo ��t��-dV�|����u7��*��˯���#��m�	��J�fR(�@�vfe�`��E�䒭��R���:H�����R�������&fhs��S��7��="���ar{�h" k�Cy �5��͜n�uV�q,��6�{X�b@��X
*,�GQ.b�Z�L/~�Μq�{Y���2�؝�[��tkJ$��Dv�
��I&���Ѕ����V��11�,?��ŒC2�]BK>�rGA���#�"��1p,.Gm����B��"vb���X;�~+��o�����y,ּ�<�Cލ�����D$�N�Vs�����޼h�]|Q�e�J@�SI�t��JC�hu�+2<	l�??fH���GE,�����#Ol�����&���t���&i燨�ې;�|�1��!��!��_9Y�6���uQ�< 0y/v!�;�Tuc�����Iĭ�	&f�c�N��gf�|B��8�����"�������q��%W]t7�����
2���J�ډ���p�v9^Ü��N�}��A�@O���&i�ېL��� �#�)�>i�oq�����tY�������
΃p�ǊY�.�N�0���k�Z�:��r��A�R� �6�L���%�?�ۆ0g��R��xb��,w
�C�}`�Y��9yq��D`HI�{bYC!�W��/R���l��7��{m���*�'I{V��
��gP&�c���Y£�ܩ�B����n���fͤ^�ARS�'w�+tz=
�pP�<=��"ǋ�`����,,K�ׂ�񝥨 Δ�|#չ����ȣ��#j{@�Jf$r��X�B�_�����1���=e����l���{:˟iv7A2ۻ�3L�3�K�1�Y�-����	{E�$���l���h��ԑ��]��SX25��e+�����&�3B��#֖H���o5,�qҏ�(K1+{�{�������q��}Ź���u���K����H54N�,	/����f�=�>̄�ʠϫ�O�`s�߈#ZO>'h]y�ܦps ;��l(����T�cˉ�T5R�F2�#o�U�p����jW/���X	�n.��Dy���-ǐ��iY~2��M;���5�R{������?~��f�3`k�]�_�[��'kQA�86�#�f�h�su��eY��⯭�䲽�ZC�Uq<�i�C�9�$ȵRc�̓/�=���_Y�K���2�l�z�6�-�eMv?�-����!����3Z"{(X��c\�O��5���h�p^+�)~��D�+BOUm�1�jT�Z[�n�4#�ǝ�B�ʽ��3���}5,z�^�4 VKߗ"�}̞�4$�R�N�$�~��f��p-W�1$����v�� �����8��N&�F��^��p?����m���݂F��s���L̩��ʙ�,�o��E�Fh��e��i{9�+o1_*��5�l=��w}����Q�A�kh�[� %��
��6'l�(\z�hj��.���w���C:%r7�(v~��p��3~&#z����:H���w���`A
�M`�f,IZd�R6�����s3@��d���Б0�>3�΃\�-�6R��u��� �'�����w��6i�+C7O��6���qpM���V|$��k��2|pKr=��gK�3��m3᫄����=�V��� fI#2:��l=������~�I��,���ݝ��[U�ѲIҏf��V0�Fs"�qlBP�����}/�S��# �I� Eh�$MY�n^BJ���nS	!9�LNg�v?\:_���4�e����UK^�m������mCR%�����>�\�?�64���G�0g#�2ષP��ox;�-�ꎢiԁ��
�õ2D~O�����xl�~ ������۬w�s��c��[�����rp��%��^T�!�����H)��ߎȞ#��
���k}��TM�ܒa:� ���.&��$��Z��E!�H#~���	�����Q�*K�LE�����4�����}�*��_����h0ʀ3�)�J����}M�b�Ԇ���۠8�����\Bv*�T^t��V}
~(42�N��TR�_�`��B�SCq���8¥]I��_e��+Շ��|�'�@R����O1D�v7==nx.>{F�,���$sB��zZ����a.,��h�Ƥ-W�~5�,%1����Ʊ筘�R{�x�$�ށcP�=Ʊ��w@�E�o�x���Yx�9�se�zNj�9p�1P��E�@v~�dh�E�/Jm�q.�S!�|��N�@64t��%�~/��P76(�f�K�sO���C1�R�o�f�hI`���%s-�`���ߌ4eY00c�����~��ڤ��g�qӺ<9��o@xW�e�Z��Wq):a��@	KX����y<0]�:7���_��ԭaN<����|g'�We�ŵ�8��)��(�ɮ�f�Nl��f}*
�M�vXѽ3���_��(p�db9�����u�V��2�AV"�
�n��2���F^0�A4q7�@�� 5�?� �����"�t��a��iV�FN�+#��}�4by���rR�n�}s��6{��}8�i�52�C�_I�3�%�H-������t���ߋ��+�2�}���{�o���K�:� ն�f5����sGT�I}ƀ��?��ރ�eB�u�͠~m1�"*�v���T݅�e����֒�G�^�K�*hSKq�{E\E��2,��3R��b00�@k��~���&a�I��XփeTu��qE���q22���Ĩ��4� /
ʓs%(��zdGXlxVHYEB    fa00    11c0$FZX�����z�����w�znI[��
�Xe�@�13�8��NM
�!��Ԏs*���b�Sr�I��DH����'�N�\�#��ɳ��DE����X	z7���f�W��	x��&i���ܡ-]�ә���Tb<�b��At�l��#F��.|Vi;��W�0��.|:�)�vq��5G�\A�R�ZQſ�Ϝ}&C�9[M�1D� 
ȝ咡����O�o㬑!���H��)]��O��M�a�T2��.�B�PmztI���i��w�W�9� �����$�5������Zk��$����O�|}���<���:$�3����thrR<��/��܍`;zK���+.���d��&��{����{�|(��,K����1F�0��m5��)EK4�ؿMNbE�c���eA�}�Us.ф�)�v��+UF{�$�ȣ$��ZG]�E���L�9 A��(#�S���P�˲����kS�N���wy:w��P�M�.&a$�.�p�Ϧ پ6D��e��T�X��jg R�ML���Ś�`r���y����,6��?2�Y5�i�h�ſ_r�)�s���!S��onJ\=�G&�i�Iýd�(T0ϧ�a�H��*?"	���P��țU'���k�`cx�?[V�a�g;",|0��l)"�L�#���Dۃ��Uv7a|sh��Ϣ������Dvg6����W�k����]w��`�=�@T3����j�s� �㓆�r�p�xD�9a�@�8����Mz5U���rB֞��V,�P{���\��=W�#�F�*[��]yv��J��a�
�m��Lk�cSBR� �qM[Z����J�W�/l��+�p�\2�%�
a�_�����ita��J���l��^$a�Х�k�%�@�'��^�~���!�A��Y�F~�j�hY�F���jU/�4��=�V��~1��8���U�V:Wj��}�.���ḏAR�x��TH�!�>�,�`ن�>
Ax��J�Y �`�-ofޡ��|m�tSu=�q�	^����9�$�H+�.'�+��N�AK�9Ug�M�~n�~����rw��y�[�$_̆�Nު%fum�;ɵ���w�{�$���g�4���G[�����ڔ��#�S��\;T�h���Uc�0��i�^�J/�M_��SՉ��F0�8�m]��NT����K��ki��]d�j��4�ẏ�H|�L����(Ӷ�� ׽ѪL +��]
͢s!� ݉�ب0���y�ZߙCm��g.��u���C�*�.�$�Cu����ovO*2��Ӵ��
9t7Eg��	!_E��({j�z��46D��'�[��)<��ŚQ��hu�f�Z��AF�ѲJp#��N.1I���j
�q��U
��-�@���c�Q)��0�Əz.no,w~-�ds������Ǆ�\�� ���s�F�*!�#?���Q���S3��дJ�ŷ$�c���f�uK7��}O����Ńr��dbT�c4k��5�{�l.^��y�L)��h@��B��p��G7}m�&d=Ӥt7A��L�5�N�8�J�v��]�`�~������5�fi��	b2��L�t�R{.��H�%�X��mIg7no� �:�)���z���Ar��<oL����vD�� ����A���HP�r�a����B��aA�`��'a��*�c��1�9��IE=�K�j�Enxt�F�L�H�4�d�R��E8ej���u��\̀	)���[�1+��7P6^T�Kp��)��MP��댴X42�aj78� hԀc�W�
�����S��i���e,qT��R1�ܒY,��C篦��f��qe��qƛ]�:_�13���l �@9����S�����*�l��&f�H@l$�e���'2ΗR�£�����Cj�Ѵ�����|zh�>A��}0��q�fG-L?�����
 �P$�)F��|G�����g���ȷ��Zy�%O@��d�,+��e՗��.�����\��^��?Qj��ԩsD�]����V��5�;h���f���gBLG3��qd�Z�k޵a���Y��i�6�TI!N�m�M|7G�t���o�֭�.�,v�t|o�x!ܦ�+?����l���:R�Hr.���]c+�W�U�AǸt��j&�m��J��r�_�)�
D����a��l���F4�co`,
�{�LN�7���@-��D�O�$Q����f�<�H�NNPK����MU�� vU�f��~L�)�MV�`�⬔����_�Oֺ���Ct���$�{����w�q
��(����&k�a���5q��Z��{ɘ��P�}��VP���L5ҼH4?�"�0;���)P�8�=��
�@)�	|�_�p�[]�g��>�H3:bb8�V~����#"ԟ!u��|��n(ۛ&G��u� �ۥ(�]�a욞<�q���.���!�7ʛno�*�f8�Hup�����(��F���*�;I���HRKCѤT��ؒM������(ObGaN7�m.;�N/����I���)��� *I�,�F" ��Q��]�����2����;h��tW�`��1���k�>�{�*����h��WI�v�6�F�r����oQٽ�O��FUm�!2�e�$�)@k3&]�U�� �T�S�ك��;��#���!d�/0�+�NVt��v2aoy�K�W]W�n�=�۷9Y�Z�M��i����6� /�
���^0S��O�E��7����"m��S �I�r����Zelu��'�{��5P�\3�'�نc��.i4)׳��Q����B��� 8"[��r�P/�D]W��\�������n*!H�>��{��П@��l,����fM���)Y/k�(.ㅸÇ�M�c:�+4���f@���o~�|�����U��3��b�(�=�];�������kTG�u1���B,Ä@�=*R#u���6�dO�^��Z�(���V1Ԛ/^zCz��1��V��,�B���{��Ɇ�.!��2���sM������.=��^r֣2c?Pڂ��z����>x�ǎ[y�}W�hOf��0sl[����T��S��Z���t��c�8��ФIAi�e����w�6a�h�:bO���(���t��D#r����:=��>���{�8��Y�����GM��S�n�~�R�K����q�^%��ND���-�%����_���N��1�6��+e���F� C%X�*��K&g�[������L���8�m�g���b����|���{7�,E�U'����_�-���I(  m�HB���T�7�{����n�y]#}2��Z����C��)%E�/�4fB���Ĳ�70��J��A*'�\	�%�`*�8W+w6C
��� �F�q���%�&�J�k�&X"d���n򑒟�6�V�G���Y��w�R�|$�;Rm���ΈF�������)�15����s�`e>^6_���=�`��i�����m�����br�Kwʠ�~��o)ETq)��3r�e�]@�7�(�ma�!�����c�T `Ծ�7!C&�U�H#���UJ�T7�/��3Zba����m�m1*3��K�ճ��|}h��c+�������F���YBN�F�ou%c��ugt䉺�,t�.�6Ӵ��d������>�Dڡ��p(�\D,aH+��+��׊�D��+�����U"�ziY��gH�z�č�r��Qo����D�����bi3y��y|��^1�&�L�f��e�3d�tXղ�5ZƔ�X=<�^dߛ�N}Fρ{�'c�9Q��'���ЛH��/��^�eg�x�t�~$o�Y��yU!�8 `*��N����}������\Y���v�)W��`�^7���~�u�|k�ϙ?���$�͸���˂B�q�9��V�����API���,�t�'0��6 ��g�`��E>�A�Ke:��:R��L0��Ӧھ����.i�s�*� �3e��,�kD���&��3��f�/UO���E��DVr���fX���+��*赆+F
��U�+�8[��V�������ڝ��uH�FټSl��<�0�'�Y�3��J�*�X�M�IS_�^�vYs�,�]ϛ�v<qӒ1m�[7��v�ҏT���4qU�Z�Iǜ�oŶ�S��b]Lm:~�p�;�7�|J�d�p�@��M.g'���/�0�����ӗ�.n8�N2S�J�� M)�g���V���h���OW�b֚BY!*�IQHk*�q����DEQ�@&}$7(H1��<tz���ߣ�F��*݇a:��鏴f~��y.n�k�P#�;ʤT~gO�':�Dfz���G��9�*��$Di��)^�����7��94���^!�-8?�4��8Q�Z4�>'�������̪����Ԥ��V���s�@z���~��oI�0?�Fְթ�{�k�%����r��/xu7G�WΗ���ׇ�#�� ۦ�6?�̱��@�f8��XlxVHYEB    fa00    2cf0�L��qO��ÿ�K��Fw��p�0^����u{�����Ѻ���H@�c�� ��=�<r�q躚��'�W;�� �H��~؊���{ϕ����p�%g�� OR��0A(�CJ����K��,!`����M��h�a�R���N�W
5|��kDZ�տ� ����H�#WϪҞ� r|K=O���%��0۷�R}��en�#ڶ�m�֔�W�۠��ĩ$��Q7��gk�$,�;z\Ehy��M$D)P�-�d�����Z������1�A�ΖH�z$�Yz-`)o<0��9�A2��� &<E���1�@2�b��q?i2�M5�oi" �B	�nŶ�(�26;�2�fԘ-7����;� �tj����b�O2@���rZ�-������HV��h`AҿW��� ����V�+�wI�|�9�i����v��扮Fnn�ə͆���{!��~w�IΤ/W2�笌+R���d���E�$��eM�����eO�����&��۽����O4��b}:2_�j`�����x�Y`���'��	�s/��Ģ'`fU�u�=����T~��M�5����k ���eِO��t{ <�����������T��骀x���t|<�ә���Yqi�?�!��?pb]ض�(�~7�L����23��a�� &��L�(7����2ˬ�6����Y�B���� ��c�61#TT�N9t�� �����n�>:� �����<_[t'O�ܟ��^�l�ꈡ����tS
�8��1����*�W���W��E�e�푝�1I��x�i(���B?�kr�v�+q���\�g+��G6\���õĔ��;��|�����M�t/j}n?��,�ʜ���Z�5����.�VV3ڍ/���.w-Ģ��ih�+\濬ܭ����fc�ag �k���Y=(�lV�ʗ}��ժ9n�h�[�pf���ݵ�*Y�~C���!�(�=�d�EI߆��Gu����4o�3=<���
3�ɚlA�ޅ��R��d\�hOp$��+(��T���E���0�`tVx��(���L���?�; Z���[�������ᶕ���.P��;���ӗ��v�L8���?n�9���и��s͉IaW��� �T��uq���F�obt���0�yu�*�?f��j9--͍xmȓ_t��\�{�b���lU[f��%{W��'�y1�Z"�rAߋb�� A!�2]z
�5<�#;Ǻ63۹�Y�	'����@wM���������YHs4�bGY�qV�gS����̞%��/&1Ӭ��lk���w�%��}�(6���C����9s�}@if����9�*~�8�~�,�FP|���k~,�����pZr�P��^��1g~"eE��>���{��6�Ц`c����7��|/K];/h�J}�g����;�$Ar.��"Amt��$r��Z:������
���j}FӤ���;��nО�;Y��|^�ZD9ms��ZfdU��)�'��r;�Tw��ݸn�c�։�H�r9��>B��	�D���VcR#c㟲m�n��c���Һo=k�5X���iA�(��S���8P�����ՅЊ!5��%��K������UO���7��ۑ����!󋳕�,_��D�dj�}���j�X�[`�q�����4�Wd
����mې�����m}� Ĩ�/���G�w��~�[���z�,�0 ���Y2��E_7�w�>��S�e���$�>t���e�jI�������4�N@TU^#ƀAC^=�aq�Mt-GI(�F,k�m��d6?�l.*�p7W@�!Z!-�k�'vX8M�Y~�wr��f�nU0�S�͟��;�m̘�?���?Z�χèF%���z�ho݈a�Q�K+�{L�E��5g�����Ɏ �_\�F	�Vv�6&�����F5h��PTZה٢��Zh~�y?��e|��8��䔑?^!ua�GQ��$�����u)�,F��`��Ώ<y�܄���(X�Ţ�l�Rya��� <����,~�[k���]B]<�߃4jQ_��I�Lv�_��uNzA�����m�[���A2���K�_��;�&��k�\��LR�_����0�l˕e��>�<���������%#��u�	��F�-?�K��{�TqP�����8�U�#-�e���0�D����"J����b1= �%ǀ�&���PU���g�olŬa�x2ۋ�xn8x�����ЍM�5�P��:2�����vOR�XD�m�Jj(ITz9&��.�����6
5AN/	zIӅ�7�o�ʚ���|�՘
eb�q������E�\4�e�*�mTJ�f�����c]&��d^ �-��=,�^�k��~?��qA�jMIp��B��n��f�f��2�ÂQ҄���+�U��W�QU{�Nk��pYE. K��k7nb����@�³t���}�𔡽E�],d
�P6�I�+=e�LP��˖���o���V6��*�Y�ɳx�#�+Cp�G/�B�:a�F>G?ZIq qPbp��Qp�����p�(kC#$�e&��-���6���P�A�ȷ�8������|yI�x{��Ag���G�}��6[\YG.f����ӥ�gM�q�`e:�I����HD��]�qC>�������G����keg4�=0�:��4¯U|`[�錉����1����.u�Ӝ�"\��>]���� ��p��	�~6d��|���@C�ӑ�t0��˱�-�ZǼ��"�`�;�R?$J��W�1�ĺ�|�!��F���;.ȼ�����d�}�?;.Y��2���LpY�p��4�##��\#G��g��]/!!U�C@����s_�t�<FR�v�a9���L�T�
�T�6��1_���l/�����Q}����P0x/��|����n�,��}l�x�eg-$�ƴ;���D<7��:���,o ?�D���J���{��\�*],����L��Z��_���s�)�����9z��g	m�X�O�u[oog9PV����B�`dd�|�T�WB�5^���*=VHf6x"|�Q��c{�~�̄o��<��S輲�K\��y{Au�`<w����F��8�<�<��ut���9;yO��0�f}j��H�X�{���/
����/׈�lj�������A��׬�x���8�]�5ݯy��t�m߇���^.q���EA��~K-��|٩��3W�P[N�JCNr�CQ�0G�y���8F���?g=�h�3�F�^,�	>C�Ω�I�ۻ'��g�A�83NwqQk�Ó�H����@~|l�ԙ(�<��A=��~�t][[cY۷������@ː��lc;����5X��c�BIKR�ýl�+y��ث��L�LR��>��AY�BL��!^#V��{� �yr4;�a�Ĥ���6�h���0�dr���_��$/6ԝ9k{�Ĥ�(OH�B�K#�O�,�� .#fT��Sk�9_����[�VB�f��E��A�KE�񥌠�4��?ɯ�H8��!�Gv�����i���uKw�/�a��G��Y: ��	�v����x>���-99'��am��}�����(Q��'�+H��Sc��D�ұ���(�}�~Wv�0�L��)5Gɩ5o>$
p�ex�X�O]��4@�୒1T�]Ip��a�}�k�}�V�c�\'X;����AL����w6���=[�1KWn��P�+��R�����ֽ��'a�zp�AۆL�o��QrF,��Ytz7���7s��XU�$L�!%��?�޽/沏h>�l:��@��95\0�+Y��𛚍Ik5
�ŰP�[2�%"�G���F�-|&J�"󸹍-$�7Q�����Qk�C�Z��֟zq���õ�����Wq&�Sx,����8CÓ�;��|��P�i4�X�r�j��-j�1�����mM��:��z=�>B|�_������uGv��� ��%����'i��Ӻ��$���!���\E��|�e$J;��-mA���0J��c5|h��(�zsM���:	������Y"�D�q�ꣿa�Y���S�U��мe�OE�1)K�n�ƞ2d���{]�%_>���DÆ}n�_F8�%��O@�t�n���0l��}姐��F��/�u(R��h�U��XnO�O���8�=�!��d��Fu
yv�i����/k!K&.����9D1����������a�kd�M����5wR;U�+��B3��"Z�6���Nm��}��������u���қ���69(#Y����,�>J�%�/��� ���Hm��2[�g�<���϶o\7�Y�r�Q��;p�ق� �,h��C���at��!�1��ЯM* ���}'�d�Y�/�g��	���b��̖��jt\�1E�ئ(%=�t������˶��be?�؇Ew�_c+Qby�����&�w�w�+��򖕅O�����06�AhT�W\�ßV!8N!��F��f�n��0[p�k�����\�1�$Ɠ���� �u��e�}r��ZR`�/[�R6Izq�`[��t�%0�!LE�Lc���޶�P#����-�`����L��t�+�f��"kNg I��~K�i�Ҟ8��,�v�/�v�C3$�"�R���	�"��Ll�	�U�	��������ƞ�C�{��������Ӽ�9�҆�z�����*h�������b`�wܱ��/;��W[�ߚ��mǯ�F�
۱�eIs����4�U|^���ۻ�Ӣo��� ���5�3�R^P�,N�=h��'x��*�9��V��Z��G�B݄�ȹ�A���l��31�G���hD��
;2Q�C[=�ËT}���JQq�S?�]L(jbAD_�m��RK�_^W~42g ��ݚ{b		{�e�]�6�l7Ŵ�DDd��/���D���d�>m\8V0���;���Q:!���9G3���c�x֟��� (a�j}�,��@���]4�*a6u����0|�l�ܶ=N�
���kYk�GW�8J�S�&]}\����<%����<�oP�?�`:D[��X^���{Yk�}i.W�J��O'G�ۢ�����R�O��5z��΃�6�Z��Q�˦:0�G�-�Ye�������Wγy��LNP���$q��hI���X���~���ޘ�����������&.������9 3r��J�^UJ%bMW�G�:CRe��?b�4�y�q�-Y�a���.��
�;����j�>T�����45��c*���\Y!b���3mT����.��|O�̽���W)cw�ٞ��Erbj�,�MP;��N:�(�<@��l��vµv�ͽ��-E�G�E^#f�4H���j�eR�ȓ@�B��8��|�qf�1s6uEX��{�-�)�&l��m�0��+�M�#l�89�f�ښ�zZ���p$��3���ݹf��ɶZB��6��/�`��
sa�5�H�,�@ݛW������c��S�|��9��o���Q�,����PB@��H���~�S�c�lєY��'�x��67H�_Vp�Xt��>ؕ2/�x�����I$D����^�'3��Z\y��1�_�Q| �f�ޏ�]�$�w�YЗNn(XI&�r`�
����`�OR� ��$�_�zg@E<�P����(������pV3���W�+��zQ_�:�����J$E���o�AW��Z��� ��V+��N
f}]���t�ҝ���x|��Q	B�a�c�=JZwq���p�jAR��k2���0v6�����^%h�ɷ�+dg�l����XR����O�qЭI��@��F�V���ɆA�.�}	���IE"���ӓ.-;d?�P�˯���	���>�jA�aBbnju1�v)��l���5������e��G�W3���8��� t�{)��d�
*O�R��N�G��嵴��v})P]��?�4���d��!?����d�1��M��AJXV�{��N�(W7B��ڬ�<��H/y/K���7��FS<c�©HH�Βӈ'�#��9�O���m����͟���c{eKo[�h'bӄ'te�m�w��o���}���T|�����%�~X�_�����_�����xi _{ 8��F$�����m��fe��^~G����T���CV0�p��� ��}��� a3���2=�o!�����u��,�����O.��X /����EG����m�tN>�! i�,�6��[s��JH^���z5�K������G�Mb=	��#j��Zxu?�.���!������"�c)f]�+G�d���	ߨ��;M5�ǂ� DZ$m�kǕ�[\�}b�����S7�ꫡ��+�:�g��Z��ke&�^��j=F�x�Й~���7�\�zP}�J�%^�s�*���F"%�-�M�����3�A�go{��;��%��2U��y���6��ޜ����3kK�fI�m5�/��87�-O)J'�.����:����'�-zͰ�R�ѡ��I�������c��h�j�-�ÈUu�B6
��u��qۄ���:/���8�ʹ10���n�~��W4-��w�1��nix�kj�&2�Gߢ����~^�YU�A��h͢��o�ny�mH�k�q�,����)��ZV��5�̡��zՑB��C<p�9��o]���T@p�ܻ�w$�k̆Z������|:��	���W]���Km)����skg]�)1�	��=�a�E�F��:��*�O|K��o���;15r8�
�.�J�~<���Ej#$NM�p�O#�2��Տ�p�}'w���b�����>������_X�հ��G����V� �<4���(��$Rn��6T�v91���þ��1"e�Zy��8J�E3T�E(ꈋls!B7��ڜ+k!���q1C�� ߩ���c�������_Ͻ]XAe�w3e�oL�zIʸ�Q�h��".Q"	�r�z'�nZ�l�΂GcL��$I|N�U�u�F^G�ڒTW��1�khT�	0.vs�O��f-���n�!��wݼ&������J��hXY�9]���a�L��&�"�PS����"o� fO?TZ|6)����<�>`������/q�!��\�b6	��I�� ���yw�,�ޕK��dam�������h:&}���b�-���x\.��u��q!踀��OWN�������	4�����j��ݹ=�X �pX��gR^@`��}���4����k�V�v[���~�����}�i�P3�#b��������Ip�Ï�>8���9�h|TE�b}g��_2���8Tvs'8T l���t�
�׭
9o��p��L"����ā�x&x${�Pf�.!:�xqPa�y�J��%�Ф��7���-#�urW3�cٵ����kvq��+��VH�-�p綸L\��=Oj����1��u�q�5��p֧�Q�_����"�����<��6�8�Ч�B���<�K*���V�i�_��^��K*���0�,B����cV���#{����C��Z��ҖGy%�r/>R��4�͊��l��ZI��<?�����ͅ*��=�e�g)O�b:X;9�}��U���E/+#on���1be����?MHk̮�;]��g�t&�Eч��n!�'1(�Ծ��h??b)8d��N����?7��i"�p���۬��$CY-Y1�J~�*�%Z���[TMH���ME*��`����X"Hq���8���C�n$�2�O�$�ի�L��s0<�z#܆@Θ<�=��t.Kep���ac�y���wT�����'��BB�)좄$�I= "��"1J�i�捔��:푨��c���1��壚-�%� P)j$)<�g�+���w� �y�.A����=go� �({L�|��ӤZ$�=i��c���d��LS8��φx8tn�Z+� @��$��TC������bʄ�	r���9l�"�U�����Ҽ6��<6	��9��
u�w~��f��ZQ�����[`h8���#zLj�8E"/Z��\�\���h����S��'�@�x:��9�s�	j���-�55�TN��R�����U6���\���x��I}�n�NS}��&q�ٮG�s�F^�����i`t��p�z!'��F~��z�Nٸ����j:Y�TL��Z����MiD�z���?�E
���K���ʕ����=a�=�}{�m����dA�k���b�D�ۜ�g��2:��#FEe�����}�Һ��8��i&���E�0��Pٮ�1=��V�\�ۡ�������|���[���XC��Y-�0`�0�U�|硑f���[���F��K2�Ԑ���w�H'�%����\�\P_�yxm�F���H<ܕ�� ~^���P�yb9=�����\El��7�5w��	9jݭlX��ޝ����
Dջ��TJ�񯨕p ��U��.���At7Xg!"uO�B0��L	S����G�z����Z��O�q�m7	���鼓k6�Uv-� ���k;Z�K`}�'k�L,��I���3%��k�의H#��j�^xZ�g��0�Qzк���^~���[���F7U�%9�>�ał���[�C�pd�_[�ل��z�;:��6]i�e�7�lswmd��1Xq�i�8rO	�zD�Ҋ��U/ !;�*�7�F�
�x��`�ꕯ����85�{���F�MRe[�a�8l�{����JD�\e������vj��+Zȋ���jb~���{13~���Zz��p4�$�;�o�,�[tZօ5�)���'j�m
�Ѩ�K֐���u��Z3�媕�=�B��'�W)�DB�a�~
�>��{y�r��J��T�)Jd^��h񨘱K��z�^}4�;|�M�e��=7ta2��+��6��L�=H'?��+���{8�?��D|䷆%~�a��$�D�ЍZ�3�/XL��\��;����Y� �v)
c9Q��Cd�Y*}��B�w\�������Mw�%c�pS�wmL��a=[Y���Ke��Z3� -�w��ס���T�w���l�'i�e	��\bX_P�a��w���6���)i�i��)�􌣺(W�6�7�Ŀr��0��&cȦ^q�9�1Ŷ��xM->��ɪ[������y	p�<��{ՙ��x��1ξ���=�S�5 �T����x�*�y� �IxEE4��
�8���:��=Rr\J���eK��C���/>o
�^~�U�NBK�p�ꎦ�P�����N}���M����Ó�VL����}D_9�����n��6g|�̀��i��d��6#���c��w*ݏ��d�>�GW-�(pzv��g����s��5��ִp�z������/fN�2��=��*j��ofL�v\�=I�rؠX�ԥ6�[g7��U�r��~�k��`Ҷ�8^�s�M�$e��;}3eJP�+��V�`�)5U����	���=��~T�U��:�d��l�:Ա{��V}��.zP�˱^Ȑ2�f�L�h{��B6Lh�G���������xr3���0Ǚbs ����P�;�Ԧ�HL}�tAm�Ŧ�î*��,���
��������ԇDF�~�x����I�h~ۻ�-�����B͡b�E�������]{{��qu#t��.$"c M��3��6�����+��l�9�?((�׌�+�Nag
��|S�շ�,��I�����g#Ekł9�h���5.'��嵀�<������!�i^�&�.����2Nyؐq�,�q�Lu��6H����>#�N����$�/�P���$w�����8F�'���sOʤ7
u�Z;r��u���ZY�w�˨�5Τ�s���DO�����w�%M��-Z���MxfH�{To��}S1<#Y����o���:y�G�x �D�I]��@��#�
���27d�諧��[�C�D��z.L"}=c���#[���-���]�0Z�o9��hbxL���K��m�4v�w�y��	���E.���l�'^�4
�AWm�a�.)�b}TU�n-��fRprٔ��٪���r��L�z����l9������L�� ����N�*������k
ԵZ�V%��Ci#��*�,�?�����zi�[�6���M�P��]<�I���~w?Z��(ŋ���{c�Z�G?JP~9�J�
m`�3����0sG�7}H��ǟ{�w`-y^���%����.T9�a+�ë�[����لk�3�
[��T�.V;���9�MF0%u(�u���%9��	��B��"x��)��OhM����a�R��`��SN�ƃ�5�$fS�G0�&fS؇8��a���}T��[�n��`:��9ݞp�~�h�5/�j��8?�%X̲���5�1�,Z�I�����E�(��sV$Z�ie��A \�5���D���]6��q�=-�XM�va9s��8��#w��7�vD��7��M.(dp ��]�BR`.�QT�v��_�|��%�=��8Э��x�_�y\N��=�;7���ĭb�2)&u���l�_o��I�ɵ.OՔ���V��]ߠk��3yla��j{]�ǛȲkcHe�n�"��6Lݹ�S?o�?{M��µ�"g��e�c�I��1y-u�2-�o���[y���[�䆕�e�OJ��c�����?K@
��)S��ꠤAA @����3�OK�8�SIn�á������9g.�~���Ls����|4�������;Ys�l�0� 泭�0�^�߮�(g)پi��Q|�Ëav��$� P�g�����K��"�$�����f$�ۧ�X�E�w ����Y{���֪M��Mt4g��p])�U�b5�
�~E�qd�&���|��R���|'B(�	٢����rX�
x����dW��sb�;m\#����:{-A��i�E
(� B�/5��7����Y�I�������>���T"���j�&V��	��m����<��!�:��齝",pǥ�:����0<lhq�>4� �ID���7|��?nipw�h2*�u.(���8zׄP�)�0�%찗�VN�!Jn�@c�a�Z�"��ܩ��U�*ӆ�}��}m�Α�� �$�ۿI��O�O��H�hh��9�?�s�H�B�y���'%HfMAN;D�9.$	��z嶃��݀��bv�4�i�BNp2}h��/��q[R&�/��	L�QO�̼W4&�"7f�JS�o��x����"�U�2��w�����?O�w�����r򜔃{\�5��P�F5�!�)�	#-u�+��K(����/7w�IEq?>�S�Q���)���3��W����#���%sv֚u.�T�z�#�k��Z�:�bmH��8�XlxVHYEB    fa00    1f60F������B��}�؇�:�������0�0�����+A�`�v�����ۘ��V��ܠA����!��N�7�u��H���6�S/n�.����D��T;�s�g�1w5��"�o�늡2tt���yGs����h�'��1+@��m�S(1ȉ��Jɼ2��#���B���,��3�kU�-�瓏�3>ͫxnJZ�pȈaSl$��1��҂���mJ���_m��z�đ�n�����XϹ��f���&Q�����D������S2�`���O�	�����^�F�m֎ӷ�C���gn]�,sz�D��vzz��b	�T�t(�z�JW�m�$(��f����s"��}����He9Qa�	���i����F3��7!de�0���4�)�Q
��"�o6�`���r5NP��Pq{�p�h>��3)����='v1�h�X�q��Ȋ]|@��e}h����8��j�����7�;r����?|�l��I�����x�bjw����Խ6�|�:���^����(������d�_�e{^��AK�a�4���$�_xL$�c�9�u򠜵�Xb��gϲ�3���� �c���6����0-����1=�By�&Q�,�^�F�����Yh��ܷ�\ā
]� q4�/q��D�����|:R��k_�o#�7s���@����@�h�kˊ3�i�"��D!�0�S�5�߈
o���.��$�.��0b ��<3=�聂dw�"��
����}|D�J%�7�QVF�n��G���w���٩��9��dL�@{cO�+s�C��5���=#ګ��_S�}�%+��k�\��G�����׼��9�
��h'����ޚ΀S�]������+xC�{��Vxr̛��Z�vnuR&wz�r������-Z���4%>/*j���e�E\h�gnw�_3�vz�ͳ�w��K�?���~��E	1C߀�s�R��y?I�ټyϢ�2M�m�gރU[��Ùv�7�}��x�@l �Y�A��'�gT�5�Pb!���W���H�f�����3&��X�^mWΒ^	�r�o>���|ڧ�m�����);^�X��.����ͼ���Ո��U]e���1dY�:�yc�G�R�E��!oh�	��I���n�lO��r��x�H1��1�Mð�������G��IB&-!��Iћ^��Hq~��{!*�26�y� �t:���
7��M��|��g�=v-�)_�!�B���%$��;}N�tfn����>U�4�X�|I�ծ�U��-�zIr��qr�'�Oæ�/,�A�J�eY%����˚�\O`�z�;�0iYZ*�X�.f��!T0��h3�b���ΧM��� [X�����#ہ�{-��=2=Iʳb��PSQ�1��T9�2�Q2s`U��(��i�2�R��N C�����J,�DR�L�̟�_���.�/�]��L9h��E;ڂu�2Z�?g����L�����R>�?�M��c[ވ1[KF�:���L����JȫY�����т��.k(��>f�}�g�SwZ��ڎa��W�ѵ���_��_۱Z�:[*�	'��^f5F��8i��g���mr�g�BJU�c��R��Hmzi������Zg8N�K���EJu%��%9�U߲!��C̆��;�ы"��Ky�z�u)�]�j�:Ы&���F�|����Ze-� ꖨjdn�ŵ �`�B�"u�kw�]�V�3
�#������d�����	��J�~#���Apc�/�]�?Dȱ}�Ab���i�r���D�Qc�pa
S�7z������Z][����\�c�����Z�_�cw¼����7?b��Ψ�����O�$M��,8����Οf�~�-N���~��M��3��x/M��A�6��`q���ǋ��'�d�/ɨm�����sh䒂��$Li��g$L��?@P�6�(V���6�Z�t(uI��F��p(�}l�)�H_�=G!-<3}͹��ᱭf�9�9	���b�m���д�D�X(�3p4u����/D�?7|fIO����x>c��P��i��ܛ�Vi�PX���U���4�/��%���H��^�ȡf���U86���ښnEen��.ǮȦՙ��׷wh���n�2ѧo����a����@/���Gs��op`���ݛqO��
��@�0"��og��+���1��_�d"�ǯ;�Ƴ��}��^w4l�����v�ݲB�9�0W��^��DN��\�Ě����(B6rP��3��q����`�bBar�7�1���g�'�> rR�k���Ş �ι?�x�D�W�lN��c�f#��9���7R9��һ��]�"� �"��թ5ur�F%���s�yl�˰��yi �R�HG��]-Pq���/
x����J
��8������(�~/�L�jl���h3]ne�'-��⤧a�_�v@˨���!�8��+( �X��/*���W���vNK��Xb�)�z+%�(M�$��������WK2+1�IA�(s"�c�[�J����Y��(#��mM�c/~�ʠzE��Hn��)An1�����P��aHEb��o�:��; @����P�J�C~�.{�@o��y���ڹ��cؿ{�ϸ<�SB8����X����~�>W\	,�P��ma�`-�`ӭP��P�ݸ<d��K��+��Ȣ#�Y��ն���@9HnSZ\�+V�O��Ӆm����Z>���Wꎥذ��5_
��:��.,&�1�I������+�����Fx���c�_mC��[^��y�*%y���!����37��hC�g���Q�;w�a��C3��d�������+	������o�B��=���j%v��V�S�k������W!�~�0`���ET�s����������Ć�%¦�Q����9�QݛqQ��i��;�zݤK@qI��9K��*��#b����� �
��
7Bh��hQ�+�3���в`�Aoxrw�&-�	|�̔F�)������tC��B{���oY� ���%�p�RJ�+�������:������?��>���dv#ךPCp����wv��~��u��	�ط%p�Bu�4,-�֙�*�&&�@o�B*_@3B�!��v0�Ըk=�!� g�����DC)��ۦ���IT�j��W�3 ��Qf���פB{N7�}?��(�#������-���3���"��:g8���wI�ᾭ����r[)�H��������l}@ g��\[R���q�Q�ٷkx4���������>`b�7��o��g[u��y2-W͵��r�}v�AKL�No��`���`�Ƴ�~��+g�6��R�F�l"��q)�=���F�Ŏ��Ӫ�;��	��nG������ж���Y��RK|�P �۫!��w�#�^�F��Y2کM�O@y�&����
 �K΅;�I�yF�/@7��ZN9���by��I2�
=�<=����(��e7��X&�e�t�e�o�a��`l��m��q���v�7����!��du�aR�9�&p��_>?>mM�)��>�;���I����@�k �;��^��;��C����:C���:Pȫ3����	 ��b�����L��Bw��'$�Z�T����F�O��l4��{�P��s��^Tm`r�,t���tx�ui~����0햡�9��%��R߰U��8Qb"�B�᯷a��,�;��m��Ǚa�Bzb��I]�ڏ�gT͡�a��c-jė��x{A,����3T��+"���2�Q�t��"Ј���y������3��sйTT��떻\�C��e!��Zq�R�M�v��-;Ǐr'�.}� �2jh�" ��q����s7�%[�P������XPagI�[$1���d;�V:D=��f��w������A���$�R�[���K �P6r��<t��?UqaVr�:��~��yu[񈽟���Ʒ;�H}V�"����Qsj0~Z��N��s"�U�Q_�g�`v�r����6��g�������sN�`�.OT�Ҍ� \�� P/G.i=��BX��l�r�h���SLxp����ش�<��&>F��Ӗ���"���w�O�O1m��=�b���#-��'x�ևD?�6���Y90Ä���ɨ�c�!��Q]��M���d�
?ct��o?�l���R� �j�ν]n�$<F�x�Oժ�����&�a��2�F�K��d-�N)"�R
�!�#�$h~.���{�@��&I�/���R*�y��hIW�����Բ�Cwdԡ�����_�䅍�Y'H]���Z���6����{?B��O�Ѳ˔2Rp<"ą�c�jELF��u�a���$NyQ��*��"8��8�`]�G�����W=��n�(*��y
�j�G���(��X�]��]h��B_� 8���Mf`���(5�~X�����4;r�{��ٽ_��w�;z/Ͽ̺�r>.��5�-��NK.U��
L��,�M[U��	��c�Y���L�-�&���x�P�qC��6�B%�ݸ-�&�rD�y#"���-�̷oK	n��T��=F �/�='�&�jܴk��j#�!h�3�|�'i�	�.P��n�l�^��=TDv���Q��5iV�7-��.�sJ�'ACۣ�Wi�jӖ>��"t�Q�	*�'>��*%@�1�ɬ�_ �]�0(dg����Zrb��z&>���iA���aj ��{.*ve�xi��7jX3���>�>?C�bW;�C��T���������-�jh�V���EA�%E=ȶ~@{�<�"S_\�h�eU�~����{��+%�z^�INF�U����5KQ�݈WID4�=NǕ�H�sB�wtAf�]�#z�f�?WPN]�	�����o�j���=LB)��R^�v�Ksh��>�'b��3/v�+�I'Rи͂N��k�A`����#\(I�i��Dc����@��թ����۠I�8�)	�.[�jT~%U��̵�p�{�zŭ��%�� ���V��0�Ł5`�MS����!���z޹��8'��D[�mW��cw�n$y���r>=p��˙�`��TO�꭛m���YlyFvc���/Z����>E����n&�<�u#�Ξ.���/ G���`�Ru���Li\ �#�����!.���q_<y ��e�#Z���O>:�4&����j���h�0���އ��ݠ��вs�W(n�����a�q�<{z�(�����;"
���un��Y��TRS��B)WpJ��?���)���y�x>��%#{ʼ�O�L|�36���`�x��b���X�Ә4r�ќ+͖J�Wz�������S�`#�/����vL��7�o���Aɒ�v����~t�!�	�!�59�'Cm�L�d���㗐`(:���<�#�^���d9���x8�O�G'>�8�q������
�����ʞ�D��Fd�N���D��3������r7�҉Ǯ3�x��O���P��:�j���5CE1�b�;�����ﲪv�1����Pԇ�HW��?�
m�&;Md)%�uYWIc�s��w���U|*C��u+�+�d�`���KW� /��7G�����t�}I�xA�&�PC%�����b<��&���b�|?�WHI��?��7��Y����&��^��4DE滠8A��[d�~d8����":�*�������QV���bS�r�5;~������F�k���R���n脻a5v�H�E,�q�!�2:����p2��g�L,��_��dF�&";C�����让�%9G�1gAFm��C��|�^�>�K1�����������J�xG�4	��X�*�T?�$��6VoNv=�b�_޷���sSu$�B�VhRc�z�?������>;ZPj-v��߅�D'w�iѕA��c�L'�cj�Y�L���]��&��.J��6`U�܊�����Ý�O�s��W5��M&<4�K�!=�B����f�}��~jbGH;P��z�0���v��8��j
�><J�Z��˷�1w��� :MѬ|�壒is���a�PS��U!�_�]])W�&�vqri�h�9*O��b�0R���c	�`r��_/��S��91���Z�-w�(������"D[�+%�Ç@����=A"�J�zˮ�N5�hc茁Ɲ=j���+IF�|~�ٔ��t���qw��b-T·��n��:��l�Fgۖb�P!-heF�-uKQw����5t<w<��U�J�9�m�[��w���K��"�o_�Dm�9˦/A �zQ�7}~��"o ��$��C��(B1�� W27���"��ԩŢUs�����]���!A��Z�`�
sm��9%�<��8�/s�y�W~�j�i��gN���?��w0�&���]���,�6��Gs/�T�D��b�X(������N��6l���Iw&{b�2i��}V'�M��c!�X}�G�����,�pӲ�4�Lj��gl�]��x�{�!�/ά�RS���lRsQ�c8r������Ȑ���<��5�v��n�������1��ԬU[�b`�
�(��k��<�J�&K��;C�1������+��x��{9s�C����h���� p�qTe��؃�j5D����#Z�!	��j�Tf>^����
�y����˲\y����j�^����8�v�?}�OmO��$�N3hh,N%!���r���Q�w=|-(��4��#�?�dt�L���K���5�O���_	����)� �G�]�0	ArY�0}QYI�֍k�F�
������	&�q��S���ԃ������s�]*J8q7X�(��bl���j���P5�?�^h�>gU8=�	6v?�I�k�I��C�G��@��)��60�r/���n{s�Omf�z���7���JT��x��HG���G�*�bWU�����#���,���(���$ŷ�{4��S�^�����}��1) �M���q��K�YN�@�G�K��pxrl�S]�gu+�cl����(�]9LY6��g�?Qi�����Jh�,���2�wU#Z���h�73�~W�O�3�F~��y�,y���⎺sHa�aԇ� s�B"�N���b��	�@���j5؃s�4_ljlRK@�$�1FS�"��PW������_LZ����׭h�H�*�fRM>wiވ�G5�٥*&a����!���n(e�N�H�f��ӕ�����*Ʌ`v3z���J&��7�37%OY[:�أ�KB8.zF�o0���koQ��R;�a��� u$T��*5n��p�5RY���T�1�D�(}����;ɬD<vx�t]�懕 ����@��即���Wk��Cˣ�t���XJ�R�u�����r�y�a�����J�f�ٲ�g��� �&�D�C��"k�����F��.�L[�fj�O�i}Qp`���i_�}Vu��ƪ?)n�+��A>�s��Ӟ�1xK��+�F���4F̐�|�=s�'(>/�`IP_E� �svq��YΈ�2�8��!�֡a3��>�X���(�b^��qf����J�(a��Gӳ.�x����NƱ�
��/[ٓbJ��[+��l�
�MMx4��lN���w�G�.���b"�0A%YY��F��,"��Hn
ˌ�M�GT8�e����$!���y! �-����}(�T�� KH�0�%��Q�NՇR?\���3��kH��h��-��V��b��9(��s�sCn�r�]�M�[ښ�=y��6PV^w�z��e��
�ѡ2�.�%���i����[����?���W��F�a%�'�~sm��?� �CӢI�,�-����^���=5� Do�-��B�Ь?�f�"H|��c۰��9���)��R/^��;�q= �>���'� �����r��E�����XlxVHYEB    cedf    1ce0�"^��9�s��{��N�=G�8���[^�2�$� ��lߟp��n(vN���a�����bƬ�4�	�C���Y�5���i��q}����'vh�'Ap�*h5�f$��ٍT��J���4A P���r�B���_����Ă��K678�22V7��׻���������	Vt��_$�΋V�SD3ݽ�B� �"�<�hh���E7����8x�董�kG�4pS��$�m]��%�m*��G��mW.*<;��L��hT����2�Qk����x���m�(�8�c��n�	p᮳̲�f�(U�k�;T��ǘl*w��Hl�S�j�;BN1?k��9�Yl6{Z�M`Y1�hڤQW�J�t�q:���N�1#p_t���t�G#�4�Ψ����E�9��]�d_�E�K��y	PW[>I6B�T9�4
_7W�Y�8�:�&,��]Txs���T������L\�j>g�R�y'��.އ(����J�¢��	�GW� 4�}��S|-��p_��`/��b����HW�8��3������c3$��ȫ��U2x/��*U3��l6@�;쯀9q`��_+�c��d�c�2�
,v�O1�Ȟ�s�_�����-Ī��+��V�x/��M��un�������DZ����:HA�VO�&�����3FQ_���z��l.�	t�x۲����������hwV�(��,tj~Qa�(hy1(e����HU�A.���'�7]�Ȩ�k$YL�)~(�b�eU����i���Y��	l섴��F�U�8�S���W@y����B��)3�T.�1��!���Ǖ{�Ȟ/o�iz���ʋ56=��,L���.�z�E�� Jrs�᭪��F��R�\�Q[���G��V4St�Z����{��b��n�䫙�㥘(� 2Io���5��U'��~����ټ����:�QV�jcx�j�a�{i��qP�R��&P�G�dk��s��%�a���`I� :�n0W�;�����Ǩ
�������6u�v�Q:Jlg5l�@�*���'�~�:�d�[��|�yq�ŠqtI�Jr�-�ڌ���f��M���-�lӂ��y�#RHtw�8 ����A�>�T�y���.O$�M�-�(���O+��{���7�=��Q�#�:R']$�A���{����x�?�[Цh4V�^<�x{B�u�Λ�s��&8	�b���y*�G�S��<>�&��\��b�
?�Kc�
 �-��I{���U�s�0Չ82r�_ĸ��B��?�Ԇ̵')��|�T���0ZǴ٥m2����;A"�R9�u�!8E��׽�G��D 0��EY�	���7�c9���C��ު������_R ��rT`#�X���0�o�'&(vK��%����j��L����%�Z	H��ӈ�@�}A7�z�|��"u�8�3�2,U �IS��c^N}�bƜ��	ŝ�v?0p���&�#�'�*u��^��$�R�-�HNW�I�[V�ݻ��*Ey��M�Ԍ_����E�c�R7��4a
��L�Fy:��8ZY��xwκ�_}}d��W�%��-���� M��8:�ي��W����#k��?^�0�{�M����X/t�$� `տ��l�Zv�� ;���w�ܜ9Y�ʗ���RH]#g��-��l��L�
�n�d���������P��:;R��}rS��I��9ze�E��0�|f��Ǚ�"s4۟�&@�Ɲ�t]m����L�nh?�x��Q������4�󾼜�!	��Ʀ� p��աD���W�oeH��bd�D����4�;����P-"/g;g`��)GBM]d�P\:T��W����C	N;ɤ�ꮟ�w����Um���Sku�Q�	���?�k�H)�!7/O�3�ZSj[�׭"�|C˺�-_�~a��O�i�E��Ք�*{�$v�ͿWk$��n��2�o	��$ִ���M�B t�>��R���$|Q��N0�,�/����� 3 ��qu���Cʃ�r�e��J�44lF _s���|��L���f��B7��0�[ �	��'�&��Fkì�j�Xp�S�K��G.��/�T-p�����m��	��~N���R_�'��$&�-�Wm��ѕ[�|J�lW���EG�������8�X֋P���Ψ��Q�\��� �u�:���M����:W��-V��T��B�''N��r���N�R�1��ʬ�z�4���4����=P`s"`��{,%��<
��j�t�s��i�0�����W1��`ZǠ��v�.���3�G���l�V��N��D�c���?�:ѕ��z1f'ή$��������ba�
�F���d����N��{�^���a��Z��W�w�4���6�I��(��%!s�)�؆A����n��嬚(����qOGB\�(�~>����* �V��8�G.3j	v+�,9:K�q�a�3�ŞOi5��HpmFuxrt.#/]"�Jx�� p���>~|�r�_�<���S%�N��u���;�_�N@�8o�G¤��d�׈܎<�n�<�'\S�!	�z!�^y��!���,��S�a�D�g	�)cͲN�\��m�8��i��"{���C�eRaJQaC���$sI�00�Yp��
�1�Et����gmna	E��+��� :S.u5��M,S֗�l	���uޣ^�?���ׄ�ʟʅ];9S�s,c^�V��RZ��tFP[�D"鞊έk���µ��Kӵ-p�0u�T��_�}��c�����Z��QK��ȼe�n��
}��Mʰ3��k�Ybw�vӮ��>�%<3��$�|*Y�L�]�KF�5Ž2�De2q����5<4�߄I��?R�M�.2"uH$P�*�Wږ�&'�'.oG�O�@<(�s��:�&�u
��s�g�a��<C����Xl<!����K�����W��*��Q�Ĳ��_TD��8�w1&�y�	�W�`h���:~q�޷��n������WL;�U�X�o&G֭X�@�E�a�K*�{	��,�t��[MXD�1UV>UH�m�zd�g�T}����>t0p.�j� q�x��[���{��$�{�a����f��)8�_���6ષ�P�M������}���`�Y7��/�������/c�~�<'St����0��}u@����:�!�*.{J���k�)6�2%i�UШ�n��_1�Ɩ�ҋ�q1�n��d��%ײ"��e�T�Q�R�0�:f/��Ϻ�~kܮ/����a�q�nV����/�̒��T�ZlRD�Ȁ�C�pg��y΢ee�'��ԗ����^�|7.z��!|.y����5������Y�C�0�7�z��� v�'����<��4�_��u��+��mO`�QU���d�K�������˻3�����dn�ƅR��#��h�f������À��ba���2��SG8�ݕ���
2�5>+D�� ���qjD:�rQ�ygQ�ê��pz��A��eg�k�F}xu� �M�Z�n�1M�B�|I&~�����+����}����g�"&K�'6rF�/fp_&?h�AI�p�Qn�R<�6��P!�w��JD������n�,��B��m}B��R�ތD��}�&L��]���I�OTS6i��.�ހF���l{�4{@���a�J�L��5u�0� E$�TC�5�
Y>6&�W�K�ci	p�P?aF*'�2(s	3DZf++k�a|�UE�}�+:]�������ÀM2NQ܇�f�e���(ձ�8vs�f��q��<�,���[�JmXw��4�1b�r[
���$�	e+wNl�'��:d���b�Ps����: ��h�����3�&>:AU�pJ� 	�S���5���ɔ�&˵2��}l���]���lb4�~���y���K�|{#'� ~@��뙸����5y�����X)��h�nG��k�0��7:��.U]�K0��p`��X�7�kT�pP�Y�E�>T�V�C��������rX��-!J|����P��Vb /���]�[?�{8subO��ý��[�μ�+FD)L��H1�Vאh?z.f��ln;��P�wݩ��=󴍘�s�\�.|/�ow{4�e����lN_Y��^��֣d�%���x���Ԝ�r@gV��W�u�^��%����)�\(Q_5yj�zO�5��Sb�?� �+��P�_yКѨ��y��~Zaٟȶ<����s��g����Z碁m?B�XfꞴ����.)<��n�(�:�C��?�����Z��G�Ii��r��� ���ZƎ�o�UɴƝ��a'������e}���f���*L�̹�DIO~EЍ�G�-����aqY���
m!\)�3^Ӟ��#�!�`~��
��v5��)�
ض��c�C\�k�o�)gꈃ�7��kv?h! a!I�V�E��CQ1&���y#/�i+s�$�vGTJ� ��&D�X�N�%�@�2���Zģ�/�B��ב�<�^=[�c�K���$��rVL8����!Q<F�q�)'�n�ol%�u�n���m*:M �e��ҭv��=���ʞ����]JŻ�
�69���rβn�=��FP�$�̷���v�85�\���X�1��ޔ�~Zf7���	+����h3�o�^���̝GfR7�^]r?���eX�R�)��|�_��L���N���3���W��lk��j�j$V����	
X���U_�5Ra��0�W?tt�T��/
�^��C��1*Bנ�Y���LS�D�|g�0��2��Pb,�iH������!iz[�躗+�T��� �\ZMi���vpb����/r�&�򝑀-�&�1��ЧLR�ʗ�"�η�GԬ֬��baGm�?��]��}U�[�T����/2@��}z������_j M�����,�EJ��4�!'���7�{T)A����U6�LX�P��!=��h��0�Z�l��?l��$�{��>���U]���? U���2ߞ;���|`]te4+��u?L���͸ɑ %����T�iZ�7������>��t$Į�(&B��#�W��(c�j��kv�T$0�g��w�⚵�=�U��|�z�Qa=? ��rT7 E����QV��f��a�-��Wic{�U�!�K��cU7ԕKV�`7�	�2[B�z�o.%�+�X���/��+U�D
i.�)�ְ`�oZ�CW�O?��,����#�d�����жq��j`D��t�NB}vg����P�Ы�ċ�f���ml����fF���:�,�|૚.�Z6��j���P���af��1���ݠ��驉9�tz����A ��d���G��E\Cr[�J�(�ݮ;4�ȃ
�����jhO�Ю�T��m��<$�C�z��ߞf�OH:�4c�B��q��Z�=�����u��6Z	�t[�f_+��F9cu��e�U9&���E����6�՞�� CЌޣ��9y�V��)C�E�/���Y,�Z�7�q�t����)�+ף)|�mCϓa�iG�(q?�M��{�sNŪ�����wT*��	U^��Q�t2rg��t�@�I��Й,�-�̀d�b1��x��b��n��	�Q�2���*2�nϯa�M,J^�F�n���&�w&���Q>�p�����oX;2ұr�d{��MG(�58Dۿ�a����!��A_"�mr}�&�6��;l��=u�]hC]?�p�skvkr�q+��R��,Na�y���}$�/�(H����� ��Vުj�Q�+�p�3h�9�k���1ƛ��[��+����	��vÈ�1;���H0?:T��ߦ�F��jb�l�Koz�YI&� Zj�r�ɖ#���:�x[���1{�!��V]��)��}!P� ���Ţ�-C�%�)�Sn���sQ�}�^"D��Gq+G ِ�J�<��v�[�������^��1�=5YZ��T��^��3P��ĒB�z�3۠Ϲ+z=O�DG��V��eʽ1�3A���Gd3rd�}w�Am�T�xR\%�`x��6�(����mu�r6�2NT���V�}�������"���4�������:&k���Or%�"-Z�����I|�S$��$�j��m�=���8`x����ͤ5<G@�LNvk����\h�u��.�X����%{�Y��>~|N��:o�Q�d+�3��
�����~����Z��yC4M�t_��.�)�f/ �k����n�dLh��+�D�����I��$n e�4�]ļ��?�FS4�D&��B�)��Hgd�O�>����7
��WNY���5ѨJ§ܳ,����H*(�h)�t�gtp�?'�f���8>���
��_���U��<���:�Z�'� ��ޯ�`0�w��]�o�����<��"Zɷ�;q�Ӳf�N:�7+=��q�&xi��Q��J; �e:����6�����o%��י����p���S������B]�8�̚�������][���$��$�@�c�� YFhf{�U���#i���X����;K�v����0�H�.-/���H�̾�͜,q_��U��I&+ć~rю�hӼ�[�3��z��YB=�w��'�uu��_Mm����YI��a�	e�x�(��G@�ct���~�j*�ħ�����ި�����#t3�8�g���A,w���3´�u�+��j�5z�Id'�GH�չ�S�A-��ޡ��M�BBpV��Ҁ�j���{��5y��$���[&I�$<Ww_�O���қnL�wY��K"@:_���_ܢά.�R���poʎ�8�����Jk�F��)�o����5d�_p8{Cu�Y�e>�W^J@�&�ؔ�I�~����ĆDr[��h�?~x��ºY#� �������Ā�V�y��%�.�Զ��y�pZ�y	�����zD��Qb¯,�6P�[���e".Gs
�$�h�j��-�t5q:�R.K { �_�������z�*'����������]�M�C�u��q�v��O��`�xq��}!S�t��x�\Dl6r�C֦�*ͬQ���h r�BB��2ހ�ͩG1��7=��yӔ1V�օ�<��vd��T��5b�����F��	�ņ�g9I�����
�~}�+�#�Ǫz��t3t�ƍu�Bj�\��ܢ+M9��'�����9j.Bz��Ή3�9�ڢ�I؆+�#�ߋM��4��ʶ�BQ��՗m��;�O�Al��o�LV�ӕH�^�(&z��~�.����CV���d���w�"��5~~��A$�lyoĹ�ׂ��lj�{�?L8����ju�J�@��6�]k<�|N�:��9����^s	�E�ID �.@)�4�u�Q�͔x� @�3p�