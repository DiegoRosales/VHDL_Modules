XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd������8���J�h!A��wLe~�&�	�z�*�p�$�	� �(�hô��KEFF�FCj�-"8����ǯ��3
�.��<�o�䮑������*��<�>щ��C�b�V�녌*{�6�6؝����5~���8+�k��Ü�x�����c�z#Q)(����e6־5���7��������_7�o�9�ۛ"�[]��8D��9F��܈��H2��ܞI���aO�l��K�Pzp'H�s��!R��� O[f;�t�U9��G�����O+��S)�#Z�7h�S?%�� H'H�=�S��2����y��O�ֲ��NO���\`�c%z!̰ȽF��*�F�$��|��f~�;���&�+����vVS>���F,��D{��0���X��H���' ��)�#�}+���N�3���j@lt�^���<�/{�y�|q��(��bԱu���K̿��R�2:{ՙF�Fu]
~�� ��oEm��Eo�"��*xC�������R=�8���xA���rN��q�Z�2�=��{ M{��wA��6��*9�������T2�uA��LT�t��C{A/a%b�P����E6n�1��I�_�����f<ۜ,#��+��·4[
�V2c�z��vx�oc�-f���f�3�)Bm�����r���,M9\�ju��-��.h{K�.b���"��i=����NÆ�aC"ϰ紳Ɇ���:V�����Wh�-���f�Y>XlxVHYEB    3d90     f60Ҋꘞ�쬋���,^�tO'/�a�Б#V���R8��I�b��1���E$'��9	�kvl[u�K�f[K&L�߶S �����f�X�ߥ��-���dPm��c�"E3]�J�#�;zO�=��6%����Q��9@dy@�6�K�)�s���]^�@�J]�|'	�"��!���p�y<�JŹ:_�L"3�<uy?��a?ʚ� F�W K?�儝2��	���4�Bg��rWb  h�=E�3�M2m�9to����t�"��h�r6�µd~��n�����$��&�.�n4�}������PǇ-�;�T8lp����o�%d�K��&�	�u��� `�9cQ��C9�[�̼��y��)��h����s~�D�ߗI��#����L�4.�.)q�G<����Cj^f(S^���}�����L���,~� H�-^�iY_B<
�/\b���m���M�;��L#��� TY��7d��Lqqt��Z�4�E:b�`Lv��nܹ+�\����V&�5x�+*� ��\���+_�ͫ7
?+�tz��
���7/�mCP�4aw(1�$�6�����u�ˁԒ�/�>�+^ ��"Dh��ۂA�q>*���p�P��kq4�̉��e�)���(D"��k�E�*!��A	Z+��^������o�bGk�#�@�z/�ُ[_���]��8�0'�����[y�i{0���D�qґ�ej�Q��jަԿ��6��򫗹
u�eҕK"�����GM5����Y���u�٬�yc�ck)j�j��Ũv/lN�7�BW2^܆�P1��k��$���ۻ/ii'�<,��~����]��`�?��!f5�C��x��&�e�4?��v!5��6�@���S&�Dv�`{ .�?|�� SS:�Jft.��l�㫲ڗM��ߢ���)^�_����(��"���ƈ�bp;m��	+<�`8�(�)A��ו�o���$m������?c�"���w@@���B����u�G{��j%�����bh*�}=.|a:w/���oS�ۆ(@c��{�P@�X-�����阘�����ǚv[@DTI��mx��A7��i�~$1��e�$���D`��_
��1ݳ}_|�=��-���ԙ��%d�\3Fx�7]�tZ�-S�b��qAk݆v1MX��v�r�摋B���-u�r��/�체O��n��Q!�.j/����׀,�����7�'��\Fo�k��o�8����kX�,��.|Ũ�.Da�%��QS���Q0��kB��k	i�#�Т�f�ݿn�r�I/��\7�XNhA������gD��	�KD���ۂ����yW�b������������P���kֆF�WaFU~9ސI�ΛlZ{�����(k��/�
LGӬ�g����R|�f���_H��	e��IyI�]D�b�����y1��#`g�N5}��fo�5Hջ�*�]��i�Fk��e.tR�Aw�;n�gj� �uQ|1L��|}����ռ����0:>�4�6: Z�ΣF�-<`�
E�;Ԟ=���~ۿI�攕U]|���>�� ��<���o�!�*���
hJE�=��L�J��#� X���&���~ā2@��Y�C�W�"�%�,��x����
���0O
~�v������Tvc�� YS�V��y5�Q�k6Ps���f��3k�)�����f�*pO�#���ŭ��`���q�����d�Q�8���ˑ�g���7L*�hF�lֺ���<�X{w+��F]��,��l�_�
zEk_��}�Q%�KKg1O�)��eNx�`�������	�1��
5!`�%��b���yZ��8bN���_�(*�6�"�8��+D���K�m�S���y^����Ay!ir�:�	xU�+�Шښ ����|��}��#U5Q�qaq��X��������;�k�1�(���J�^�#�9B�o�`X�`K$3�\�#D.�7U4�26�,4!nr܆Y��q��Fu3jg-ؕ#�����D�>ř{0��)�W�n��	S�ImV1^_~`	^�4��l��y>%��)�>�Q�^�#^��o��m�i�`XE~$���-s��G"������i�[�*��-)i��6hFpQM��j<�9o�qOk�ָ"�gl���Ӡ�0V�p�X��>�e�$�Q3FhK�n�	��wzPE���0@�飁M|`y����D�wۦ��l/ȵy{u���}�
rk8:*HB���
h?Ԭ�QW�;����j z�W=+<!!�����a�THc7��@AЎw<� J���i�tvI�cC��p(��š�w�A�������b/��S�Q�e�u��h/G�<a��X�6�C۾�����Ó�&��+�	�y!���c����Z�S�fKDC��,���.�O`>��)�_LG9�a�˗U莅@N�����F,�?���+k�
R��)��h�~ �MQ��p��4n[�,΋@��0�,A����e,K�i���jp��B3.��-|���Lg�tf5��8���'�Q�e*��D!��E���4~V����7p}��<QB��q<s�Ww"M����=t2�c
�d=^�uO�HV�����"Gܷס���AI��ߵU�H�א��~'O��P퉴!o�hb��p[��*S�Gvх+ݹt�V��;b��=J㹇,Ғ��b���8�g�ED�QQ���LtI�f�7ޱ�ի�������v�P���Z"H�|N��ȹ1�	�Y{V!0\1gxS�����5�����AE�LG�K���𾒱���Ro$C�V-��Wg&@o���a����6*�ƦJ;�= �/5�x�6/2{1�3$N��8̐�;=��݉2)o`wF�+�g���x��xm�EY�����D���\�W?����8]��zt���[m䰪@�h�D���w���~̴?@�m�`��寬f�[��z��Y��)���mDki�hL���u{�� ٔ�G�qg=�I^�T�c{!�݈v�7{x��kiޜ��`���Zj��I�<�>Hx�q�sH�?BsC�}�5O=!��P�Z|�ಭ�%ש���Sɾ����D���A��R.�0	��$�4�n�I�4���a�6O����.��Jm�vS��t+.�At!���1D^/�Áz�Ԟl4Gl_�-<iH�3J�~�\�$n�^�_�ވ��
�qu4��N�8�����]V�7֊3�K�;�"��Y@㏌�����ݧ��}���=�~ʫ�t�gi�ɒD�ۡ+�J�I�����)'!
&�ְ,�K>�����;ЦF�pp�h��L#$��yH�׬i�\YV(�κ�^�,�P�.�=y}�U�L�"Ǎ��![�I�H\Q�9 ��
���ֆ=rD0��)�Zj�$���MAWp�gİ��DX�
O�����W�BQ֕�b(�yEm�-Z��ze�ǉ��W�J?c�ϡ�u4���x�EC2��2�%�O�U�仼g�o���u�������n��D��[�&۪�bt�%�
��T���]#r2��^U����$�#��.�
�)�׸&��C��R�jB�J��Z5���\^G25��Ad.)�C+��� �<�;_��U�em禄q�"�<��N#�d����ʒ���}E��E���!/2@47O��?a8�\ �<h0�k� ����A�=�==��/.�H�*�aeM1}���Bm~��RO0�_���B�KZSa�[�+U0�zW�\͑j8��S��&N�,�R�KPs��c��V�y����*�k.�2�����[�GIl�m������ra�K��\�g��E �Ey!�gE<�OP[�9 h8,���IHrF1nW�3芡ZMR�_;��[���