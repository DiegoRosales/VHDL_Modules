XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��ҹ���>����5Bi�?���[�Jdp�@�\�D�o,¹��
�[B �0�y�KK,lS;6��;I,�$�a�H�o�v��{�n:EҰ��x�_��vX[U���D�c�Z���s���0�Epr�� ma��u(^nvWf��='͓4i��<O��j?8;��[r�=	����<pӡ�n���Y�OU���-J]ޢ^�\AxD�i��\�^�d��وO$4W�D½ ��LP�4�k{�z(j��r�=��tk���ݴ�PH&��Z�E6�/��Z�v?^öZ�*�n�1�ڏ.�����#:�[��9��9��V�F���;1?tA�y�,Ma~Lp�v�܉T8�d�E�r�W�JQX���[�d5���,�5����7�F4�B���Ha4��J����m�`���WX��E�"���Qg�v�r�*�)f3�>^>x
{�T)��9qaY�J@�;%7Ě�:�R�p����5b
&�#~���f�|zc���@�|�h.@�|�2�re{�6��ݵ[���A2��.���%. R���x�w�����i�h<ְc�W��-�G���N���uV��c�8���U#���Hᄊ�*y�S���l{nVq_�B�������8��s�ǔK��t�m+���qd�d����XE�3� F� k и'to����_Ի�m?�vil�!�����/� ����'�($�R��P�K��K�7Tt�9,����{o�oN�u��d��X�ֳ�O�ia���R���VR�{�|2`:XlxVHYEB    2bbe     c70x ;��|��F���@�8d~;,�J���m�-z����v?�<��#z �K��E=};��	��ş��߀";��0����0
=����S�)&1�� �C�� �!_�;`�f4S���k�h��Iv�r��e=��G��V�^4{}[ y�ב�Ե��|���,��n��1��R�F:
�!���,�;	�"�oi2'�:�u�Z����(���;��T.{8��� :<��R
��a�&��� �,�%�P��R��К;Vy�ÚÉ�+%�~�g�+��|5�����)�yU�YRo
�CU�x�� ���&��+�̷e-s�|N��}����||P��A$�z;�A���'
�N{�L�c�u�zX=߀�.��ەce�	"S�=L�B���������Q��1� e�'�zd���k�_�В	��Z�����> �
q0L�CWT p��g�t�[�����������?J�ў���Oiw�/��QD��H
P��u�3S�C��u�|���U�99w������6���/p��h��������q�&E � �u���[��2��Җ��7[f;t���m�r���ɚ�>�gXjW�kCU��z�ǉ9(u �A`žH'إg�w}��Y��wT�b=�WH���`?>��hV��hb�I(1���H-+ï��}dީB���M>�� �q�H0���,ēɡl�$������[B�Va�B��/Ҋ�%��"�n9ĝy[G�9=	~�\��n��`I�ϹAS2�`q@�\�#�@��<)�b3�Ik�z!T�fAQ<;���u�+��su�b��||���ˠ�˱�*����q������2��-��!�G^�R<��M e=�,�3��^�M���b1�m����y�� ,�� �E���RP3%	��ib� ���]�Mr@]�6��^[�_���|�)
Qw��L4��q�'��"�a��-���Sv�,������-vh�5߯Xc�t�)�������S���;� �lǁ1u�|�*l�FCp���>G�}���D�2 �w��#k�,Lǆ�G�]r�2�fwXq�:�,�����[=�(R�H��Z�6�\
����c$[`Y/@nuw_����ͼ^�=k�O�eY�yWM�F`O�f��d���-��Cm<�;u��,������3A�u?xZ�2��� �z���4+el��U�S�v(���E���+1]��l���	�d;xِ�(}�����&2<�R=�[�ۍ��J)��_}hY6:�i�iB�Ö ��3uj�h����ۣ�?��{'ow@:+k���F�Ɂ"�vX|�*�u�8{�#t�RH��G1�&`�����*�Kf��#��Wk���L��i��4i\����!i
tc�����"蕂�ʫ�J�&�@j�6�)%�%:]�^3�Ȱ��_ꍣ�8�̔�[� �r!��h0�<&SӞ�XՏS�r�[�)���>�[D~K%0!F�l�q�!��A�o���h[�u��Z�J����)�� ���E8�.U�$�^���D�w[�[��?����W�g�B5,��ݻJ���%^�7�b��(���7T�'�2���U��5�� ��r!��r���Q�h��:��@:���Bl��_X�lH������:���衔ZM�	���*�k�#�q*d8 �)�7���7���;�$(T������/!@ܵt/���Ng�aKww��[J�?)F�u$Gq��scʼ� )���ǘ6���J����Scm��˱L}��@s�=#i�J(6_�0�-�ؽq(O!�ZӇ���2��o1�Zҹ��ld�����$g���䩚�M3ĚZ����������+��/v�_�[!o�$S�t/i[���#���k10!T�'.f�Ɋ��$�1me��Q]�U����.ϓ��ᆴҒ`;��^��ImhӐ�.�`zj]w�,��<2|�j���b#QH5`���0
��YZ�Ķ�:����]�9�v�4�{��x��	�ZF��e�Sp�~��`uEa�o�gU4el!zg����C�&�w�߼~i2�-�?���Sb��$���̤ ��-����V!�j��nu������P�Z���QQ�cp Q��a��`��B���xɽ���k�}��:�Ɵ]@{&��*�3��3�QcM�Lj���+�\�MU��۟O�w�rN��1XHa�a�����b���N��G�����</η��Gs3f�;#yX=�%��N,C�s�{	q�ۧ��(F��o;7����+E�������A���6KRoY����_]�gSs��&��?J�:h�f�b��^Sj�,7�tx��͓��b������B�fQe��q����\g��8�^��@�������;�ߨs�{2)��uC����	�q�� �ֵ�
%iB)P��٫!Ǖ�9ψP����A�Z�dg��<�R#�*۲��1�Cp�V��:������-�$1�	�*л�3�Y+S�&�<줙�5�դ+\�R<Υ�&�\�k_����4�K�(�=I�����z��V��-8��~����Q��u�T��L����32��<9�A�_1���s��?��gW��,�Vd�p�M�Ws۝���@8�Ed���>�p+�Mv Q���bS�bqHg=�
���2�d��k����#�Ly(+����8V�#6zX[���_ ����/F�J#�Kw�	�t��%�®} �z�	7����E�s���˹>��	�.��F���]����X��$��2����d��z��ٸ����΢���HFˠz�+/���tTp�m �PNxV��a�=օ�&���JĐ���W����#���������Fmy�&
�A^ �RQ˛j��)����oj��F~���
UCt��4�u�Ϝ�t���׍�4��>w֧W���u�&T��0YU~��i���p܀���9�_����Q�h{�����U��Kj��{�K��<��Tu��羣��l�-nxhx�톜�(�7��C�%-�O A���$�uԹ�Q�S��bi��$T�a�}5�^g4��y \
7&�V�_�*�����?T���J1AP���p +\}_��h�Q.%* �"�H��OM��t