XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��7��	 +s�6)*`��uE*E !�|,up_Z��p�-,�e�!�;��Iz��J�f2Ac0�5A/�F@�fĀy\0��啱5R�$��qdO�a�8�d��\�p�6Z�*�zŪ�ՓO�v; >�(�+}��</{rٝ�U�/�[Z��@>��[��1ʲ�lTҴ�( ��X_߶��֊�a�\�N�;�4��i�Ao6g<�� u0|h������a���5���Ga
�4!�g�4��Ď}l)��뀔q�M[\̰���q��j���]�
[�/����ֳe�UB�fs�
��z��!�9,;�j����9sBh�_�2'�öC�7L��;'p̸\���Ӵ�v���v:���hj�����e�#�}څ�ݴz��:/���>��5IYm� �6r��);	e,�_�����cp)_�i�9�������k�(�Ϧw��+�̈�f"?�J�#�1�d|���/�:�K<��7��$��$}��0�{��.�NLG��|A5�}c���Q`K纤�;�#��x�[�Й!6�	��1�w6�C���0���+���r1;�&p5 d�du��	gS�q'��Ep��ݻ�6�E�l-'	�H
��Ӷ����K�K�O�?��� MM�zſ!�e޴'{�O��� ���]��Jl*sW}vq�a�)]����x#~B֑u1Y�%�G,-��QJP0��)�8���k�34Eh��Fm��I�5�� ��b�B�T�3�M"��!��!�x���um�XlxVHYEB     872     290я$��L�ʹ� �f"q�ה�F�%,ͣ�x��N9ٲ��|
��PȚ���-�1�O�Rvr�EB��B��q���y<�8ōt`��"����.�ր�4�!K��"��`�N 0�6h�Us�q��}�ׅ156W�ͪuo#�)��<`?��lf	���'��k���:�-�D��R�;���T�����&�yU�@��HvO���2ź�����0|���3\��מ�O������c�VZ�rUq�K��im�̎�h9�ҝ��,ZeI����L��-�.鐸�XP�|�|���@�^�'G�(�(x��u�	'@�c�?j`��EL�l�m��hr��C����#� ���mbգ��'�^}�f6���|�1h��=��O��A��1)��!��I���T�7죋��yK��kq�/!yj�;��pw��݄f���bdP/�#XY2��x#9�'Fm5�F��0�a�Q[�{��J�z�/�(<��nY嘟Q�h����%�n'Vq�yrm򤸞>�*��5���kv�6�9:���=媊�A�_���}Cpw&����Z;�I@/!����9�����V�� rw`p�"F��EU���*
�:�ʙ�k�����ȳ��o�ސv�!���iz�孂j�N